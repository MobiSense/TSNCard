`timescale 1ns / 1ps

module ab_traffic_exp_switch_tb;
    
    parameter TB_MODE = "DEMO";
    // parameter FRAME_LENGTH = 1514;
    parameter FRAME_LENGTH = 1400;

    // `define FRAME_TYP [8*62+62+62+8*4+4+4+8*4+4+4+1:1]
    `define FRAME_TYP [8*1516+1516+1516+8*4+4+4+8*4+4+4+1:1]

    tri_mode_ethernet_mac_0_max_frame_typ frame0();
    tri_mode_ethernet_mac_0_max_frame_typ frame1();
    tri_mode_ethernet_mac_0_max_frame_typ frame2();
    tri_mode_ethernet_mac_0_max_frame_typ frame3();

    tri_mode_ethernet_mac_0_max_frame_typ rx_stimulus_working_frame_0();
    tri_mode_ethernet_mac_0_max_frame_typ rx_stimulus_working_frame_1();
    tri_mode_ethernet_mac_0_max_frame_typ rx_stimulus_working_frame_2();
    tri_mode_ethernet_mac_0_max_frame_typ rx_stimulus_working_frame_3();
    tri_mode_ethernet_mac_0_max_frame_typ tx_monitor_working_frame_0();
    tri_mode_ethernet_mac_0_max_frame_typ tx_monitor_working_frame_1();
    tri_mode_ethernet_mac_0_max_frame_typ tx_monitor_working_frame_2();
    tri_mode_ethernet_mac_0_max_frame_typ tx_monitor_working_frame_3();

    integer i_stimulus; // loop variable
    integer i_monitor; // loop variable
    integer payload_length;

    //----------------------------------------------------------------------------
    // Stimulus - Frame data
    //----------------------------------------------------------------------------
    // The following constant holds the stimulus for the testbench. It is
    // an ordered array of frames, with frame 0 the first to be injected
    // into the core transmit interface by the testbench.
    //----------------------------------------------------------------------------
    initial
    begin
        //-----------
        // Frame 0
        //-----------
        frame0.data[0]  = 8'h00;  frame0.valid[0]  = 1'b1;  frame0.error[0]  = 1'b0; // Destination Address (03)
        frame0.data[1]  = 8'h00;  frame0.valid[1]  = 1'b1;  frame0.error[1]  = 1'b0;
        frame0.data[2]  = 8'h00;  frame0.valid[2]  = 1'b1;  frame0.error[2]  = 1'b0;
        frame0.data[3]  = 8'h00;  frame0.valid[3]  = 1'b1;  frame0.error[3]  = 1'b0;
        frame0.data[4]  = 8'h00;  frame0.valid[4]  = 1'b1;  frame0.error[4]  = 1'b0;
        frame0.data[5]  = 8'h03;  frame0.valid[5]  = 1'b1;  frame0.error[5]  = 1'b0;
        frame0.data[6]  = 8'h00;  frame0.valid[6]  = 1'b1;  frame0.error[6]  = 1'b0; // Source Address  (01)
        frame0.data[7]  = 8'h00;  frame0.valid[7]  = 1'b1;  frame0.error[7]  = 1'b0;
        frame0.data[8]  = 8'h00;  frame0.valid[8]  = 1'b1;  frame0.error[8]  = 1'b0;
        frame0.data[9]  = 8'h00;  frame0.valid[9]  = 1'b1;  frame0.error[9]  = 1'b0;
        frame0.data[10] = 8'h00;  frame0.valid[10] = 1'b1;  frame0.error[10] = 1'b0;
        frame0.data[11] = 8'h01;  frame0.valid[11] = 1'b1;  frame0.error[11] = 1'b0;
        frame0.data[12] = 8'h81;  frame0.valid[12] = 1'b1;  frame0.error[12] = 1'b0;
        frame0.data[13] = 8'h00;  frame0.valid[13] = 1'b1;  frame0.error[13] = 1'b0; // Length/Type = Length = 1500

        frame0.data[  14] = 8'h00; frame0.valid[  14] = 1'b1; frame0.error[  14] = 1'b0;frame0.data[  15] = 8'h01; frame0.valid[  15] = 1'b1; frame0.error[  15] = 1'b0;frame0.data[  16] = 8'h02; frame0.valid[  16] = 1'b1; frame0.error[  16] = 1'b0;frame0.data[  17] = 8'h03; frame0.valid[  17] = 1'b1; frame0.error[  17] = 1'b0;frame0.data[  18] = 8'h04; frame0.valid[  18] = 1'b1; frame0.error[  18] = 1'b0;frame0.data[  19] = 8'h05; frame0.valid[  19] = 1'b1; frame0.error[  19] = 1'b0;frame0.data[  20] = 8'h06; frame0.valid[  20] = 1'b1; frame0.error[  20] = 1'b0;frame0.data[  21] = 8'h07; frame0.valid[  21] = 1'b1; frame0.error[  21] = 1'b0;frame0.data[  22] = 8'h08; frame0.valid[  22] = 1'b1; frame0.error[  22] = 1'b0;frame0.data[  23] = 8'h09; frame0.valid[  23] = 1'b1; frame0.error[  23] = 1'b0;frame0.data[  24] = 8'h0A; frame0.valid[  24] = 1'b1; frame0.error[  24] = 1'b0;frame0.data[  25] = 8'h0B; frame0.valid[  25] = 1'b1; frame0.error[  25] = 1'b0;frame0.data[  26] = 8'h0C; frame0.valid[  26] = 1'b1; frame0.error[  26] = 1'b0;frame0.data[  27] = 8'h0D; frame0.valid[  27] = 1'b1; frame0.error[  27] = 1'b0;frame0.data[  28] = 8'h0E; frame0.valid[  28] = 1'b1; frame0.error[  28] = 1'b0;frame0.data[  29] = 8'h0F; frame0.valid[  29] = 1'b1; frame0.error[  29] = 1'b0;
        frame0.data[  30] = 8'h10; frame0.valid[  30] = 1'b1; frame0.error[  30] = 1'b0;frame0.data[  31] = 8'h11; frame0.valid[  31] = 1'b1; frame0.error[  31] = 1'b0;frame0.data[  32] = 8'h12; frame0.valid[  32] = 1'b1; frame0.error[  32] = 1'b0;frame0.data[  33] = 8'h13; frame0.valid[  33] = 1'b1; frame0.error[  33] = 1'b0;frame0.data[  34] = 8'h14; frame0.valid[  34] = 1'b1; frame0.error[  34] = 1'b0;frame0.data[  35] = 8'h15; frame0.valid[  35] = 1'b1; frame0.error[  35] = 1'b0;frame0.data[  36] = 8'h16; frame0.valid[  36] = 1'b1; frame0.error[  36] = 1'b0;frame0.data[  37] = 8'h17; frame0.valid[  37] = 1'b1; frame0.error[  37] = 1'b0;frame0.data[  38] = 8'h18; frame0.valid[  38] = 1'b1; frame0.error[  38] = 1'b0;frame0.data[  39] = 8'h19; frame0.valid[  39] = 1'b1; frame0.error[  39] = 1'b0;frame0.data[  40] = 8'h1A; frame0.valid[  40] = 1'b1; frame0.error[  40] = 1'b0;frame0.data[  41] = 8'h1B; frame0.valid[  41] = 1'b1; frame0.error[  41] = 1'b0;frame0.data[  42] = 8'h1C; frame0.valid[  42] = 1'b1; frame0.error[  42] = 1'b0;frame0.data[  43] = 8'h1D; frame0.valid[  43] = 1'b1; frame0.error[  43] = 1'b0;frame0.data[  44] = 8'h1E; frame0.valid[  44] = 1'b1; frame0.error[  44] = 1'b0;frame0.data[  45] = 8'h1F; frame0.valid[  45] = 1'b1; frame0.error[  45] = 1'b0;
        frame0.data[  46] = 8'h20; frame0.valid[  46] = 1'b1; frame0.error[  46] = 1'b0;frame0.data[  47] = 8'h21; frame0.valid[  47] = 1'b1; frame0.error[  47] = 1'b0;frame0.data[  48] = 8'h22; frame0.valid[  48] = 1'b1; frame0.error[  48] = 1'b0;frame0.data[  49] = 8'h23; frame0.valid[  49] = 1'b1; frame0.error[  49] = 1'b0;frame0.data[  50] = 8'h24; frame0.valid[  50] = 1'b1; frame0.error[  50] = 1'b0;frame0.data[  51] = 8'h25; frame0.valid[  51] = 1'b1; frame0.error[  51] = 1'b0;frame0.data[  52] = 8'h26; frame0.valid[  52] = 1'b1; frame0.error[  52] = 1'b0;frame0.data[  53] = 8'h27; frame0.valid[  53] = 1'b1; frame0.error[  53] = 1'b0;frame0.data[  54] = 8'h28; frame0.valid[  54] = 1'b1; frame0.error[  54] = 1'b0;frame0.data[  55] = 8'h29; frame0.valid[  55] = 1'b1; frame0.error[  55] = 1'b0;frame0.data[  56] = 8'h2A; frame0.valid[  56] = 1'b1; frame0.error[  56] = 1'b0;frame0.data[  57] = 8'h2B; frame0.valid[  57] = 1'b1; frame0.error[  57] = 1'b0;frame0.data[  58] = 8'h2C; frame0.valid[  58] = 1'b1; frame0.error[  58] = 1'b0;frame0.data[  59] = 8'h2D; frame0.valid[  59] = 1'b1; frame0.error[  59] = 1'b0;frame0.data[  60] = 8'h2E; frame0.valid[  60] = 1'b1; frame0.error[  60] = 1'b0;frame0.data[  61] = 8'h2F; frame0.valid[  61] = 1'b1; frame0.error[  61] = 1'b0;
        frame0.data[  62] = 8'h30; frame0.valid[  62] = 1'b1; frame0.error[  62] = 1'b0;frame0.data[  63] = 8'h31; frame0.valid[  63] = 1'b1; frame0.error[  63] = 1'b0;frame0.data[  64] = 8'h32; frame0.valid[  64] = 1'b1; frame0.error[  64] = 1'b0;frame0.data[  65] = 8'h33; frame0.valid[  65] = 1'b1; frame0.error[  65] = 1'b0;frame0.data[  66] = 8'h34; frame0.valid[  66] = 1'b1; frame0.error[  66] = 1'b0;frame0.data[  67] = 8'h35; frame0.valid[  67] = 1'b1; frame0.error[  67] = 1'b0;frame0.data[  68] = 8'h36; frame0.valid[  68] = 1'b1; frame0.error[  68] = 1'b0;frame0.data[  69] = 8'h37; frame0.valid[  69] = 1'b1; frame0.error[  69] = 1'b0;frame0.data[  70] = 8'h38; frame0.valid[  70] = 1'b1; frame0.error[  70] = 1'b0;frame0.data[  71] = 8'h39; frame0.valid[  71] = 1'b1; frame0.error[  71] = 1'b0;frame0.data[  72] = 8'h3A; frame0.valid[  72] = 1'b1; frame0.error[  72] = 1'b0;frame0.data[  73] = 8'h3B; frame0.valid[  73] = 1'b1; frame0.error[  73] = 1'b0;frame0.data[  74] = 8'h3C; frame0.valid[  74] = 1'b1; frame0.error[  74] = 1'b0;frame0.data[  75] = 8'h3D; frame0.valid[  75] = 1'b1; frame0.error[  75] = 1'b0;frame0.data[  76] = 8'h3E; frame0.valid[  76] = 1'b1; frame0.error[  76] = 1'b0;frame0.data[  77] = 8'h3F; frame0.valid[  77] = 1'b1; frame0.error[  77] = 1'b0;
        frame0.data[  78] = 8'h40; frame0.valid[  78] = 1'b1; frame0.error[  78] = 1'b0;frame0.data[  79] = 8'h41; frame0.valid[  79] = 1'b1; frame0.error[  79] = 1'b0;frame0.data[  80] = 8'h42; frame0.valid[  80] = 1'b1; frame0.error[  80] = 1'b0;frame0.data[  81] = 8'h43; frame0.valid[  81] = 1'b1; frame0.error[  81] = 1'b0;frame0.data[  82] = 8'h44; frame0.valid[  82] = 1'b1; frame0.error[  82] = 1'b0;frame0.data[  83] = 8'h45; frame0.valid[  83] = 1'b1; frame0.error[  83] = 1'b0;frame0.data[  84] = 8'h46; frame0.valid[  84] = 1'b1; frame0.error[  84] = 1'b0;frame0.data[  85] = 8'h47; frame0.valid[  85] = 1'b1; frame0.error[  85] = 1'b0;frame0.data[  86] = 8'h48; frame0.valid[  86] = 1'b1; frame0.error[  86] = 1'b0;frame0.data[  87] = 8'h49; frame0.valid[  87] = 1'b1; frame0.error[  87] = 1'b0;frame0.data[  88] = 8'h4A; frame0.valid[  88] = 1'b1; frame0.error[  88] = 1'b0;frame0.data[  89] = 8'h4B; frame0.valid[  89] = 1'b1; frame0.error[  89] = 1'b0;frame0.data[  90] = 8'h4C; frame0.valid[  90] = 1'b1; frame0.error[  90] = 1'b0;frame0.data[  91] = 8'h4D; frame0.valid[  91] = 1'b1; frame0.error[  91] = 1'b0;frame0.data[  92] = 8'h4E; frame0.valid[  92] = 1'b1; frame0.error[  92] = 1'b0;frame0.data[  93] = 8'h4F; frame0.valid[  93] = 1'b1; frame0.error[  93] = 1'b0;
        frame0.data[  94] = 8'h50; frame0.valid[  94] = 1'b1; frame0.error[  94] = 1'b0;frame0.data[  95] = 8'h51; frame0.valid[  95] = 1'b1; frame0.error[  95] = 1'b0;frame0.data[  96] = 8'h52; frame0.valid[  96] = 1'b1; frame0.error[  96] = 1'b0;frame0.data[  97] = 8'h53; frame0.valid[  97] = 1'b1; frame0.error[  97] = 1'b0;frame0.data[  98] = 8'h54; frame0.valid[  98] = 1'b1; frame0.error[  98] = 1'b0;frame0.data[  99] = 8'h55; frame0.valid[  99] = 1'b1; frame0.error[  99] = 1'b0;frame0.data[ 100] = 8'h56; frame0.valid[ 100] = 1'b1; frame0.error[ 100] = 1'b0;frame0.data[ 101] = 8'h57; frame0.valid[ 101] = 1'b1; frame0.error[ 101] = 1'b0;frame0.data[ 102] = 8'h58; frame0.valid[ 102] = 1'b1; frame0.error[ 102] = 1'b0;frame0.data[ 103] = 8'h59; frame0.valid[ 103] = 1'b1; frame0.error[ 103] = 1'b0;frame0.data[ 104] = 8'h5A; frame0.valid[ 104] = 1'b1; frame0.error[ 104] = 1'b0;frame0.data[ 105] = 8'h5B; frame0.valid[ 105] = 1'b1; frame0.error[ 105] = 1'b0;frame0.data[ 106] = 8'h5C; frame0.valid[ 106] = 1'b1; frame0.error[ 106] = 1'b0;frame0.data[ 107] = 8'h5D; frame0.valid[ 107] = 1'b1; frame0.error[ 107] = 1'b0;frame0.data[ 108] = 8'h5E; frame0.valid[ 108] = 1'b1; frame0.error[ 108] = 1'b0;frame0.data[ 109] = 8'h5F; frame0.valid[ 109] = 1'b1; frame0.error[ 109] = 1'b0;
        frame0.data[ 110] = 8'h60; frame0.valid[ 110] = 1'b1; frame0.error[ 110] = 1'b0;frame0.data[ 111] = 8'h61; frame0.valid[ 111] = 1'b1; frame0.error[ 111] = 1'b0;frame0.data[ 112] = 8'h62; frame0.valid[ 112] = 1'b1; frame0.error[ 112] = 1'b0;frame0.data[ 113] = 8'h63; frame0.valid[ 113] = 1'b1; frame0.error[ 113] = 1'b0;frame0.data[ 114] = 8'h64; frame0.valid[ 114] = 1'b1; frame0.error[ 114] = 1'b0;frame0.data[ 115] = 8'h65; frame0.valid[ 115] = 1'b1; frame0.error[ 115] = 1'b0;frame0.data[ 116] = 8'h66; frame0.valid[ 116] = 1'b1; frame0.error[ 116] = 1'b0;frame0.data[ 117] = 8'h67; frame0.valid[ 117] = 1'b1; frame0.error[ 117] = 1'b0;frame0.data[ 118] = 8'h68; frame0.valid[ 118] = 1'b1; frame0.error[ 118] = 1'b0;frame0.data[ 119] = 8'h69; frame0.valid[ 119] = 1'b1; frame0.error[ 119] = 1'b0;frame0.data[ 120] = 8'h6A; frame0.valid[ 120] = 1'b1; frame0.error[ 120] = 1'b0;frame0.data[ 121] = 8'h6B; frame0.valid[ 121] = 1'b1; frame0.error[ 121] = 1'b0;frame0.data[ 122] = 8'h6C; frame0.valid[ 122] = 1'b1; frame0.error[ 122] = 1'b0;frame0.data[ 123] = 8'h6D; frame0.valid[ 123] = 1'b1; frame0.error[ 123] = 1'b0;frame0.data[ 124] = 8'h6E; frame0.valid[ 124] = 1'b1; frame0.error[ 124] = 1'b0;frame0.data[ 125] = 8'h6F; frame0.valid[ 125] = 1'b1; frame0.error[ 125] = 1'b0;
        frame0.data[ 126] = 8'h70; frame0.valid[ 126] = 1'b1; frame0.error[ 126] = 1'b0;frame0.data[ 127] = 8'h71; frame0.valid[ 127] = 1'b1; frame0.error[ 127] = 1'b0;frame0.data[ 128] = 8'h72; frame0.valid[ 128] = 1'b1; frame0.error[ 128] = 1'b0;frame0.data[ 129] = 8'h73; frame0.valid[ 129] = 1'b1; frame0.error[ 129] = 1'b0;frame0.data[ 130] = 8'h74; frame0.valid[ 130] = 1'b1; frame0.error[ 130] = 1'b0;frame0.data[ 131] = 8'h75; frame0.valid[ 131] = 1'b1; frame0.error[ 131] = 1'b0;frame0.data[ 132] = 8'h76; frame0.valid[ 132] = 1'b1; frame0.error[ 132] = 1'b0;frame0.data[ 133] = 8'h77; frame0.valid[ 133] = 1'b1; frame0.error[ 133] = 1'b0;frame0.data[ 134] = 8'h78; frame0.valid[ 134] = 1'b1; frame0.error[ 134] = 1'b0;frame0.data[ 135] = 8'h79; frame0.valid[ 135] = 1'b1; frame0.error[ 135] = 1'b0;frame0.data[ 136] = 8'h7A; frame0.valid[ 136] = 1'b1; frame0.error[ 136] = 1'b0;frame0.data[ 137] = 8'h7B; frame0.valid[ 137] = 1'b1; frame0.error[ 137] = 1'b0;frame0.data[ 138] = 8'h7C; frame0.valid[ 138] = 1'b1; frame0.error[ 138] = 1'b0;frame0.data[ 139] = 8'h7D; frame0.valid[ 139] = 1'b1; frame0.error[ 139] = 1'b0;frame0.data[ 140] = 8'h7E; frame0.valid[ 140] = 1'b1; frame0.error[ 140] = 1'b0;frame0.data[ 141] = 8'h7F; frame0.valid[ 141] = 1'b1; frame0.error[ 141] = 1'b0;
        frame0.data[ 142] = 8'h80; frame0.valid[ 142] = 1'b1; frame0.error[ 142] = 1'b0;frame0.data[ 143] = 8'h81; frame0.valid[ 143] = 1'b1; frame0.error[ 143] = 1'b0;frame0.data[ 144] = 8'h82; frame0.valid[ 144] = 1'b1; frame0.error[ 144] = 1'b0;frame0.data[ 145] = 8'h83; frame0.valid[ 145] = 1'b1; frame0.error[ 145] = 1'b0;frame0.data[ 146] = 8'h84; frame0.valid[ 146] = 1'b1; frame0.error[ 146] = 1'b0;frame0.data[ 147] = 8'h85; frame0.valid[ 147] = 1'b1; frame0.error[ 147] = 1'b0;frame0.data[ 148] = 8'h86; frame0.valid[ 148] = 1'b1; frame0.error[ 148] = 1'b0;frame0.data[ 149] = 8'h87; frame0.valid[ 149] = 1'b1; frame0.error[ 149] = 1'b0;frame0.data[ 150] = 8'h88; frame0.valid[ 150] = 1'b1; frame0.error[ 150] = 1'b0;frame0.data[ 151] = 8'h89; frame0.valid[ 151] = 1'b1; frame0.error[ 151] = 1'b0;frame0.data[ 152] = 8'h8A; frame0.valid[ 152] = 1'b1; frame0.error[ 152] = 1'b0;frame0.data[ 153] = 8'h8B; frame0.valid[ 153] = 1'b1; frame0.error[ 153] = 1'b0;frame0.data[ 154] = 8'h8C; frame0.valid[ 154] = 1'b1; frame0.error[ 154] = 1'b0;frame0.data[ 155] = 8'h8D; frame0.valid[ 155] = 1'b1; frame0.error[ 155] = 1'b0;frame0.data[ 156] = 8'h8E; frame0.valid[ 156] = 1'b1; frame0.error[ 156] = 1'b0;frame0.data[ 157] = 8'h8F; frame0.valid[ 157] = 1'b1; frame0.error[ 157] = 1'b0;
        frame0.data[ 158] = 8'h90; frame0.valid[ 158] = 1'b1; frame0.error[ 158] = 1'b0;frame0.data[ 159] = 8'h91; frame0.valid[ 159] = 1'b1; frame0.error[ 159] = 1'b0;frame0.data[ 160] = 8'h92; frame0.valid[ 160] = 1'b1; frame0.error[ 160] = 1'b0;frame0.data[ 161] = 8'h93; frame0.valid[ 161] = 1'b1; frame0.error[ 161] = 1'b0;frame0.data[ 162] = 8'h94; frame0.valid[ 162] = 1'b1; frame0.error[ 162] = 1'b0;frame0.data[ 163] = 8'h95; frame0.valid[ 163] = 1'b1; frame0.error[ 163] = 1'b0;frame0.data[ 164] = 8'h96; frame0.valid[ 164] = 1'b1; frame0.error[ 164] = 1'b0;frame0.data[ 165] = 8'h97; frame0.valid[ 165] = 1'b1; frame0.error[ 165] = 1'b0;frame0.data[ 166] = 8'h98; frame0.valid[ 166] = 1'b1; frame0.error[ 166] = 1'b0;frame0.data[ 167] = 8'h99; frame0.valid[ 167] = 1'b1; frame0.error[ 167] = 1'b0;frame0.data[ 168] = 8'h9A; frame0.valid[ 168] = 1'b1; frame0.error[ 168] = 1'b0;frame0.data[ 169] = 8'h9B; frame0.valid[ 169] = 1'b1; frame0.error[ 169] = 1'b0;frame0.data[ 170] = 8'h9C; frame0.valid[ 170] = 1'b1; frame0.error[ 170] = 1'b0;frame0.data[ 171] = 8'h9D; frame0.valid[ 171] = 1'b1; frame0.error[ 171] = 1'b0;frame0.data[ 172] = 8'h9E; frame0.valid[ 172] = 1'b1; frame0.error[ 172] = 1'b0;frame0.data[ 173] = 8'h9F; frame0.valid[ 173] = 1'b1; frame0.error[ 173] = 1'b0;
        frame0.data[ 174] = 8'hA0; frame0.valid[ 174] = 1'b1; frame0.error[ 174] = 1'b0;frame0.data[ 175] = 8'hA1; frame0.valid[ 175] = 1'b1; frame0.error[ 175] = 1'b0;frame0.data[ 176] = 8'hA2; frame0.valid[ 176] = 1'b1; frame0.error[ 176] = 1'b0;frame0.data[ 177] = 8'hA3; frame0.valid[ 177] = 1'b1; frame0.error[ 177] = 1'b0;frame0.data[ 178] = 8'hA4; frame0.valid[ 178] = 1'b1; frame0.error[ 178] = 1'b0;frame0.data[ 179] = 8'hA5; frame0.valid[ 179] = 1'b1; frame0.error[ 179] = 1'b0;frame0.data[ 180] = 8'hA6; frame0.valid[ 180] = 1'b1; frame0.error[ 180] = 1'b0;frame0.data[ 181] = 8'hA7; frame0.valid[ 181] = 1'b1; frame0.error[ 181] = 1'b0;frame0.data[ 182] = 8'hA8; frame0.valid[ 182] = 1'b1; frame0.error[ 182] = 1'b0;frame0.data[ 183] = 8'hA9; frame0.valid[ 183] = 1'b1; frame0.error[ 183] = 1'b0;frame0.data[ 184] = 8'hAA; frame0.valid[ 184] = 1'b1; frame0.error[ 184] = 1'b0;frame0.data[ 185] = 8'hAB; frame0.valid[ 185] = 1'b1; frame0.error[ 185] = 1'b0;frame0.data[ 186] = 8'hAC; frame0.valid[ 186] = 1'b1; frame0.error[ 186] = 1'b0;frame0.data[ 187] = 8'hAD; frame0.valid[ 187] = 1'b1; frame0.error[ 187] = 1'b0;frame0.data[ 188] = 8'hAE; frame0.valid[ 188] = 1'b1; frame0.error[ 188] = 1'b0;frame0.data[ 189] = 8'hAF; frame0.valid[ 189] = 1'b1; frame0.error[ 189] = 1'b0;
        frame0.data[ 190] = 8'hB0; frame0.valid[ 190] = 1'b1; frame0.error[ 190] = 1'b0;frame0.data[ 191] = 8'hB1; frame0.valid[ 191] = 1'b1; frame0.error[ 191] = 1'b0;frame0.data[ 192] = 8'hB2; frame0.valid[ 192] = 1'b1; frame0.error[ 192] = 1'b0;frame0.data[ 193] = 8'hB3; frame0.valid[ 193] = 1'b1; frame0.error[ 193] = 1'b0;frame0.data[ 194] = 8'hB4; frame0.valid[ 194] = 1'b1; frame0.error[ 194] = 1'b0;frame0.data[ 195] = 8'hB5; frame0.valid[ 195] = 1'b1; frame0.error[ 195] = 1'b0;frame0.data[ 196] = 8'hB6; frame0.valid[ 196] = 1'b1; frame0.error[ 196] = 1'b0;frame0.data[ 197] = 8'hB7; frame0.valid[ 197] = 1'b1; frame0.error[ 197] = 1'b0;frame0.data[ 198] = 8'hB8; frame0.valid[ 198] = 1'b1; frame0.error[ 198] = 1'b0;frame0.data[ 199] = 8'hB9; frame0.valid[ 199] = 1'b1; frame0.error[ 199] = 1'b0;frame0.data[ 200] = 8'hBA; frame0.valid[ 200] = 1'b1; frame0.error[ 200] = 1'b0;frame0.data[ 201] = 8'hBB; frame0.valid[ 201] = 1'b1; frame0.error[ 201] = 1'b0;frame0.data[ 202] = 8'hBC; frame0.valid[ 202] = 1'b1; frame0.error[ 202] = 1'b0;frame0.data[ 203] = 8'hBD; frame0.valid[ 203] = 1'b1; frame0.error[ 203] = 1'b0;frame0.data[ 204] = 8'hBE; frame0.valid[ 204] = 1'b1; frame0.error[ 204] = 1'b0;frame0.data[ 205] = 8'hBF; frame0.valid[ 205] = 1'b1; frame0.error[ 205] = 1'b0;
        frame0.data[ 206] = 8'hC0; frame0.valid[ 206] = 1'b1; frame0.error[ 206] = 1'b0;frame0.data[ 207] = 8'hC1; frame0.valid[ 207] = 1'b1; frame0.error[ 207] = 1'b0;frame0.data[ 208] = 8'hC2; frame0.valid[ 208] = 1'b1; frame0.error[ 208] = 1'b0;frame0.data[ 209] = 8'hC3; frame0.valid[ 209] = 1'b1; frame0.error[ 209] = 1'b0;frame0.data[ 210] = 8'hC4; frame0.valid[ 210] = 1'b1; frame0.error[ 210] = 1'b0;frame0.data[ 211] = 8'hC5; frame0.valid[ 211] = 1'b1; frame0.error[ 211] = 1'b0;frame0.data[ 212] = 8'hC6; frame0.valid[ 212] = 1'b1; frame0.error[ 212] = 1'b0;frame0.data[ 213] = 8'hC7; frame0.valid[ 213] = 1'b1; frame0.error[ 213] = 1'b0;frame0.data[ 214] = 8'hC8; frame0.valid[ 214] = 1'b1; frame0.error[ 214] = 1'b0;frame0.data[ 215] = 8'hC9; frame0.valid[ 215] = 1'b1; frame0.error[ 215] = 1'b0;frame0.data[ 216] = 8'hCA; frame0.valid[ 216] = 1'b1; frame0.error[ 216] = 1'b0;frame0.data[ 217] = 8'hCB; frame0.valid[ 217] = 1'b1; frame0.error[ 217] = 1'b0;frame0.data[ 218] = 8'hCC; frame0.valid[ 218] = 1'b1; frame0.error[ 218] = 1'b0;frame0.data[ 219] = 8'hCD; frame0.valid[ 219] = 1'b1; frame0.error[ 219] = 1'b0;frame0.data[ 220] = 8'hCE; frame0.valid[ 220] = 1'b1; frame0.error[ 220] = 1'b0;frame0.data[ 221] = 8'hCF; frame0.valid[ 221] = 1'b1; frame0.error[ 221] = 1'b0;
        frame0.data[ 222] = 8'hD0; frame0.valid[ 222] = 1'b1; frame0.error[ 222] = 1'b0;frame0.data[ 223] = 8'hD1; frame0.valid[ 223] = 1'b1; frame0.error[ 223] = 1'b0;frame0.data[ 224] = 8'hD2; frame0.valid[ 224] = 1'b1; frame0.error[ 224] = 1'b0;frame0.data[ 225] = 8'hD3; frame0.valid[ 225] = 1'b1; frame0.error[ 225] = 1'b0;frame0.data[ 226] = 8'hD4; frame0.valid[ 226] = 1'b1; frame0.error[ 226] = 1'b0;frame0.data[ 227] = 8'hD5; frame0.valid[ 227] = 1'b1; frame0.error[ 227] = 1'b0;frame0.data[ 228] = 8'hD6; frame0.valid[ 228] = 1'b1; frame0.error[ 228] = 1'b0;frame0.data[ 229] = 8'hD7; frame0.valid[ 229] = 1'b1; frame0.error[ 229] = 1'b0;frame0.data[ 230] = 8'hD8; frame0.valid[ 230] = 1'b1; frame0.error[ 230] = 1'b0;frame0.data[ 231] = 8'hD9; frame0.valid[ 231] = 1'b1; frame0.error[ 231] = 1'b0;frame0.data[ 232] = 8'hDA; frame0.valid[ 232] = 1'b1; frame0.error[ 232] = 1'b0;frame0.data[ 233] = 8'hDB; frame0.valid[ 233] = 1'b1; frame0.error[ 233] = 1'b0;frame0.data[ 234] = 8'hDC; frame0.valid[ 234] = 1'b1; frame0.error[ 234] = 1'b0;frame0.data[ 235] = 8'hDD; frame0.valid[ 235] = 1'b1; frame0.error[ 235] = 1'b0;frame0.data[ 236] = 8'hDE; frame0.valid[ 236] = 1'b1; frame0.error[ 236] = 1'b0;frame0.data[ 237] = 8'hDF; frame0.valid[ 237] = 1'b1; frame0.error[ 237] = 1'b0;
        frame0.data[ 238] = 8'hE0; frame0.valid[ 238] = 1'b1; frame0.error[ 238] = 1'b0;frame0.data[ 239] = 8'hE1; frame0.valid[ 239] = 1'b1; frame0.error[ 239] = 1'b0;frame0.data[ 240] = 8'hE2; frame0.valid[ 240] = 1'b1; frame0.error[ 240] = 1'b0;frame0.data[ 241] = 8'hE3; frame0.valid[ 241] = 1'b1; frame0.error[ 241] = 1'b0;frame0.data[ 242] = 8'hE4; frame0.valid[ 242] = 1'b1; frame0.error[ 242] = 1'b0;frame0.data[ 243] = 8'hE5; frame0.valid[ 243] = 1'b1; frame0.error[ 243] = 1'b0;frame0.data[ 244] = 8'hE6; frame0.valid[ 244] = 1'b1; frame0.error[ 244] = 1'b0;frame0.data[ 245] = 8'hE7; frame0.valid[ 245] = 1'b1; frame0.error[ 245] = 1'b0;frame0.data[ 246] = 8'hE8; frame0.valid[ 246] = 1'b1; frame0.error[ 246] = 1'b0;frame0.data[ 247] = 8'hE9; frame0.valid[ 247] = 1'b1; frame0.error[ 247] = 1'b0;frame0.data[ 248] = 8'hEA; frame0.valid[ 248] = 1'b1; frame0.error[ 248] = 1'b0;frame0.data[ 249] = 8'hEB; frame0.valid[ 249] = 1'b1; frame0.error[ 249] = 1'b0;frame0.data[ 250] = 8'hEC; frame0.valid[ 250] = 1'b1; frame0.error[ 250] = 1'b0;frame0.data[ 251] = 8'hED; frame0.valid[ 251] = 1'b1; frame0.error[ 251] = 1'b0;frame0.data[ 252] = 8'hEE; frame0.valid[ 252] = 1'b1; frame0.error[ 252] = 1'b0;frame0.data[ 253] = 8'hEF; frame0.valid[ 253] = 1'b1; frame0.error[ 253] = 1'b0;
        frame0.data[ 254] = 8'hF0; frame0.valid[ 254] = 1'b1; frame0.error[ 254] = 1'b0;frame0.data[ 255] = 8'hF1; frame0.valid[ 255] = 1'b1; frame0.error[ 255] = 1'b0;frame0.data[ 256] = 8'hF2; frame0.valid[ 256] = 1'b1; frame0.error[ 256] = 1'b0;frame0.data[ 257] = 8'hF3; frame0.valid[ 257] = 1'b1; frame0.error[ 257] = 1'b0;frame0.data[ 258] = 8'hF4; frame0.valid[ 258] = 1'b1; frame0.error[ 258] = 1'b0;frame0.data[ 259] = 8'hF5; frame0.valid[ 259] = 1'b1; frame0.error[ 259] = 1'b0;frame0.data[ 260] = 8'hF6; frame0.valid[ 260] = 1'b1; frame0.error[ 260] = 1'b0;frame0.data[ 261] = 8'hF7; frame0.valid[ 261] = 1'b1; frame0.error[ 261] = 1'b0;frame0.data[ 262] = 8'hF8; frame0.valid[ 262] = 1'b1; frame0.error[ 262] = 1'b0;frame0.data[ 263] = 8'hF9; frame0.valid[ 263] = 1'b1; frame0.error[ 263] = 1'b0;frame0.data[ 264] = 8'hFA; frame0.valid[ 264] = 1'b1; frame0.error[ 264] = 1'b0;frame0.data[ 265] = 8'hFB; frame0.valid[ 265] = 1'b1; frame0.error[ 265] = 1'b0;frame0.data[ 266] = 8'hFC; frame0.valid[ 266] = 1'b1; frame0.error[ 266] = 1'b0;frame0.data[ 267] = 8'hFD; frame0.valid[ 267] = 1'b1; frame0.error[ 267] = 1'b0;frame0.data[ 268] = 8'hFE; frame0.valid[ 268] = 1'b1; frame0.error[ 268] = 1'b0;frame0.data[ 269] = 8'h00; frame0.valid[ 269] = 1'b1; frame0.error[ 269] = 1'b0;
        frame0.data[ 270] = 8'h01; frame0.valid[ 270] = 1'b1; frame0.error[ 270] = 1'b0;frame0.data[ 271] = 8'h02; frame0.valid[ 271] = 1'b1; frame0.error[ 271] = 1'b0;frame0.data[ 272] = 8'h03; frame0.valid[ 272] = 1'b1; frame0.error[ 272] = 1'b0;frame0.data[ 273] = 8'h04; frame0.valid[ 273] = 1'b1; frame0.error[ 273] = 1'b0;frame0.data[ 274] = 8'h05; frame0.valid[ 274] = 1'b1; frame0.error[ 274] = 1'b0;frame0.data[ 275] = 8'h06; frame0.valid[ 275] = 1'b1; frame0.error[ 275] = 1'b0;frame0.data[ 276] = 8'h07; frame0.valid[ 276] = 1'b1; frame0.error[ 276] = 1'b0;frame0.data[ 277] = 8'h08; frame0.valid[ 277] = 1'b1; frame0.error[ 277] = 1'b0;frame0.data[ 278] = 8'h09; frame0.valid[ 278] = 1'b1; frame0.error[ 278] = 1'b0;frame0.data[ 279] = 8'h0A; frame0.valid[ 279] = 1'b1; frame0.error[ 279] = 1'b0;frame0.data[ 280] = 8'h0B; frame0.valid[ 280] = 1'b1; frame0.error[ 280] = 1'b0;frame0.data[ 281] = 8'h0C; frame0.valid[ 281] = 1'b1; frame0.error[ 281] = 1'b0;frame0.data[ 282] = 8'h0D; frame0.valid[ 282] = 1'b1; frame0.error[ 282] = 1'b0;frame0.data[ 283] = 8'h0E; frame0.valid[ 283] = 1'b1; frame0.error[ 283] = 1'b0;frame0.data[ 284] = 8'h0F; frame0.valid[ 284] = 1'b1; frame0.error[ 284] = 1'b0;frame0.data[ 285] = 8'h10; frame0.valid[ 285] = 1'b1; frame0.error[ 285] = 1'b0;
        frame0.data[ 286] = 8'h11; frame0.valid[ 286] = 1'b1; frame0.error[ 286] = 1'b0;frame0.data[ 287] = 8'h12; frame0.valid[ 287] = 1'b1; frame0.error[ 287] = 1'b0;frame0.data[ 288] = 8'h13; frame0.valid[ 288] = 1'b1; frame0.error[ 288] = 1'b0;frame0.data[ 289] = 8'h14; frame0.valid[ 289] = 1'b1; frame0.error[ 289] = 1'b0;frame0.data[ 290] = 8'h15; frame0.valid[ 290] = 1'b1; frame0.error[ 290] = 1'b0;frame0.data[ 291] = 8'h16; frame0.valid[ 291] = 1'b1; frame0.error[ 291] = 1'b0;frame0.data[ 292] = 8'h17; frame0.valid[ 292] = 1'b1; frame0.error[ 292] = 1'b0;frame0.data[ 293] = 8'h18; frame0.valid[ 293] = 1'b1; frame0.error[ 293] = 1'b0;frame0.data[ 294] = 8'h19; frame0.valid[ 294] = 1'b1; frame0.error[ 294] = 1'b0;frame0.data[ 295] = 8'h1A; frame0.valid[ 295] = 1'b1; frame0.error[ 295] = 1'b0;frame0.data[ 296] = 8'h1B; frame0.valid[ 296] = 1'b1; frame0.error[ 296] = 1'b0;frame0.data[ 297] = 8'h1C; frame0.valid[ 297] = 1'b1; frame0.error[ 297] = 1'b0;frame0.data[ 298] = 8'h1D; frame0.valid[ 298] = 1'b1; frame0.error[ 298] = 1'b0;frame0.data[ 299] = 8'h1E; frame0.valid[ 299] = 1'b1; frame0.error[ 299] = 1'b0;frame0.data[ 300] = 8'h1F; frame0.valid[ 300] = 1'b1; frame0.error[ 300] = 1'b0;frame0.data[ 301] = 8'h20; frame0.valid[ 301] = 1'b1; frame0.error[ 301] = 1'b0;
        frame0.data[ 302] = 8'h21; frame0.valid[ 302] = 1'b1; frame0.error[ 302] = 1'b0;frame0.data[ 303] = 8'h22; frame0.valid[ 303] = 1'b1; frame0.error[ 303] = 1'b0;frame0.data[ 304] = 8'h23; frame0.valid[ 304] = 1'b1; frame0.error[ 304] = 1'b0;frame0.data[ 305] = 8'h24; frame0.valid[ 305] = 1'b1; frame0.error[ 305] = 1'b0;frame0.data[ 306] = 8'h25; frame0.valid[ 306] = 1'b1; frame0.error[ 306] = 1'b0;frame0.data[ 307] = 8'h26; frame0.valid[ 307] = 1'b1; frame0.error[ 307] = 1'b0;frame0.data[ 308] = 8'h27; frame0.valid[ 308] = 1'b1; frame0.error[ 308] = 1'b0;frame0.data[ 309] = 8'h28; frame0.valid[ 309] = 1'b1; frame0.error[ 309] = 1'b0;frame0.data[ 310] = 8'h29; frame0.valid[ 310] = 1'b1; frame0.error[ 310] = 1'b0;frame0.data[ 311] = 8'h2A; frame0.valid[ 311] = 1'b1; frame0.error[ 311] = 1'b0;frame0.data[ 312] = 8'h2B; frame0.valid[ 312] = 1'b1; frame0.error[ 312] = 1'b0;frame0.data[ 313] = 8'h2C; frame0.valid[ 313] = 1'b1; frame0.error[ 313] = 1'b0;frame0.data[ 314] = 8'h2D; frame0.valid[ 314] = 1'b1; frame0.error[ 314] = 1'b0;frame0.data[ 315] = 8'h2E; frame0.valid[ 315] = 1'b1; frame0.error[ 315] = 1'b0;frame0.data[ 316] = 8'h2F; frame0.valid[ 316] = 1'b1; frame0.error[ 316] = 1'b0;frame0.data[ 317] = 8'h30; frame0.valid[ 317] = 1'b1; frame0.error[ 317] = 1'b0;
        frame0.data[ 318] = 8'h31; frame0.valid[ 318] = 1'b1; frame0.error[ 318] = 1'b0;frame0.data[ 319] = 8'h32; frame0.valid[ 319] = 1'b1; frame0.error[ 319] = 1'b0;frame0.data[ 320] = 8'h33; frame0.valid[ 320] = 1'b1; frame0.error[ 320] = 1'b0;frame0.data[ 321] = 8'h34; frame0.valid[ 321] = 1'b1; frame0.error[ 321] = 1'b0;frame0.data[ 322] = 8'h35; frame0.valid[ 322] = 1'b1; frame0.error[ 322] = 1'b0;frame0.data[ 323] = 8'h36; frame0.valid[ 323] = 1'b1; frame0.error[ 323] = 1'b0;frame0.data[ 324] = 8'h37; frame0.valid[ 324] = 1'b1; frame0.error[ 324] = 1'b0;frame0.data[ 325] = 8'h38; frame0.valid[ 325] = 1'b1; frame0.error[ 325] = 1'b0;frame0.data[ 326] = 8'h39; frame0.valid[ 326] = 1'b1; frame0.error[ 326] = 1'b0;frame0.data[ 327] = 8'h3A; frame0.valid[ 327] = 1'b1; frame0.error[ 327] = 1'b0;frame0.data[ 328] = 8'h3B; frame0.valid[ 328] = 1'b1; frame0.error[ 328] = 1'b0;frame0.data[ 329] = 8'h3C; frame0.valid[ 329] = 1'b1; frame0.error[ 329] = 1'b0;frame0.data[ 330] = 8'h3D; frame0.valid[ 330] = 1'b1; frame0.error[ 330] = 1'b0;frame0.data[ 331] = 8'h3E; frame0.valid[ 331] = 1'b1; frame0.error[ 331] = 1'b0;frame0.data[ 332] = 8'h3F; frame0.valid[ 332] = 1'b1; frame0.error[ 332] = 1'b0;frame0.data[ 333] = 8'h40; frame0.valid[ 333] = 1'b1; frame0.error[ 333] = 1'b0;
        frame0.data[ 334] = 8'h41; frame0.valid[ 334] = 1'b1; frame0.error[ 334] = 1'b0;frame0.data[ 335] = 8'h42; frame0.valid[ 335] = 1'b1; frame0.error[ 335] = 1'b0;frame0.data[ 336] = 8'h43; frame0.valid[ 336] = 1'b1; frame0.error[ 336] = 1'b0;frame0.data[ 337] = 8'h44; frame0.valid[ 337] = 1'b1; frame0.error[ 337] = 1'b0;frame0.data[ 338] = 8'h45; frame0.valid[ 338] = 1'b1; frame0.error[ 338] = 1'b0;frame0.data[ 339] = 8'h46; frame0.valid[ 339] = 1'b1; frame0.error[ 339] = 1'b0;frame0.data[ 340] = 8'h47; frame0.valid[ 340] = 1'b1; frame0.error[ 340] = 1'b0;frame0.data[ 341] = 8'h48; frame0.valid[ 341] = 1'b1; frame0.error[ 341] = 1'b0;frame0.data[ 342] = 8'h49; frame0.valid[ 342] = 1'b1; frame0.error[ 342] = 1'b0;frame0.data[ 343] = 8'h4A; frame0.valid[ 343] = 1'b1; frame0.error[ 343] = 1'b0;frame0.data[ 344] = 8'h4B; frame0.valid[ 344] = 1'b1; frame0.error[ 344] = 1'b0;frame0.data[ 345] = 8'h4C; frame0.valid[ 345] = 1'b1; frame0.error[ 345] = 1'b0;frame0.data[ 346] = 8'h4D; frame0.valid[ 346] = 1'b1; frame0.error[ 346] = 1'b0;frame0.data[ 347] = 8'h4E; frame0.valid[ 347] = 1'b1; frame0.error[ 347] = 1'b0;frame0.data[ 348] = 8'h4F; frame0.valid[ 348] = 1'b1; frame0.error[ 348] = 1'b0;frame0.data[ 349] = 8'h50; frame0.valid[ 349] = 1'b1; frame0.error[ 349] = 1'b0;
        frame0.data[ 350] = 8'h51; frame0.valid[ 350] = 1'b1; frame0.error[ 350] = 1'b0;frame0.data[ 351] = 8'h52; frame0.valid[ 351] = 1'b1; frame0.error[ 351] = 1'b0;frame0.data[ 352] = 8'h53; frame0.valid[ 352] = 1'b1; frame0.error[ 352] = 1'b0;frame0.data[ 353] = 8'h54; frame0.valid[ 353] = 1'b1; frame0.error[ 353] = 1'b0;frame0.data[ 354] = 8'h55; frame0.valid[ 354] = 1'b1; frame0.error[ 354] = 1'b0;frame0.data[ 355] = 8'h56; frame0.valid[ 355] = 1'b1; frame0.error[ 355] = 1'b0;frame0.data[ 356] = 8'h57; frame0.valid[ 356] = 1'b1; frame0.error[ 356] = 1'b0;frame0.data[ 357] = 8'h58; frame0.valid[ 357] = 1'b1; frame0.error[ 357] = 1'b0;frame0.data[ 358] = 8'h59; frame0.valid[ 358] = 1'b1; frame0.error[ 358] = 1'b0;frame0.data[ 359] = 8'h5A; frame0.valid[ 359] = 1'b1; frame0.error[ 359] = 1'b0;frame0.data[ 360] = 8'h5B; frame0.valid[ 360] = 1'b1; frame0.error[ 360] = 1'b0;frame0.data[ 361] = 8'h5C; frame0.valid[ 361] = 1'b1; frame0.error[ 361] = 1'b0;frame0.data[ 362] = 8'h5D; frame0.valid[ 362] = 1'b1; frame0.error[ 362] = 1'b0;frame0.data[ 363] = 8'h5E; frame0.valid[ 363] = 1'b1; frame0.error[ 363] = 1'b0;frame0.data[ 364] = 8'h5F; frame0.valid[ 364] = 1'b1; frame0.error[ 364] = 1'b0;frame0.data[ 365] = 8'h60; frame0.valid[ 365] = 1'b1; frame0.error[ 365] = 1'b0;
        frame0.data[ 366] = 8'h61; frame0.valid[ 366] = 1'b1; frame0.error[ 366] = 1'b0;frame0.data[ 367] = 8'h62; frame0.valid[ 367] = 1'b1; frame0.error[ 367] = 1'b0;frame0.data[ 368] = 8'h63; frame0.valid[ 368] = 1'b1; frame0.error[ 368] = 1'b0;frame0.data[ 369] = 8'h64; frame0.valid[ 369] = 1'b1; frame0.error[ 369] = 1'b0;frame0.data[ 370] = 8'h65; frame0.valid[ 370] = 1'b1; frame0.error[ 370] = 1'b0;frame0.data[ 371] = 8'h66; frame0.valid[ 371] = 1'b1; frame0.error[ 371] = 1'b0;frame0.data[ 372] = 8'h67; frame0.valid[ 372] = 1'b1; frame0.error[ 372] = 1'b0;frame0.data[ 373] = 8'h68; frame0.valid[ 373] = 1'b1; frame0.error[ 373] = 1'b0;frame0.data[ 374] = 8'h69; frame0.valid[ 374] = 1'b1; frame0.error[ 374] = 1'b0;frame0.data[ 375] = 8'h6A; frame0.valid[ 375] = 1'b1; frame0.error[ 375] = 1'b0;frame0.data[ 376] = 8'h6B; frame0.valid[ 376] = 1'b1; frame0.error[ 376] = 1'b0;frame0.data[ 377] = 8'h6C; frame0.valid[ 377] = 1'b1; frame0.error[ 377] = 1'b0;frame0.data[ 378] = 8'h6D; frame0.valid[ 378] = 1'b1; frame0.error[ 378] = 1'b0;frame0.data[ 379] = 8'h6E; frame0.valid[ 379] = 1'b1; frame0.error[ 379] = 1'b0;frame0.data[ 380] = 8'h6F; frame0.valid[ 380] = 1'b1; frame0.error[ 380] = 1'b0;frame0.data[ 381] = 8'h70; frame0.valid[ 381] = 1'b1; frame0.error[ 381] = 1'b0;
        frame0.data[ 382] = 8'h71; frame0.valid[ 382] = 1'b1; frame0.error[ 382] = 1'b0;frame0.data[ 383] = 8'h72; frame0.valid[ 383] = 1'b1; frame0.error[ 383] = 1'b0;frame0.data[ 384] = 8'h73; frame0.valid[ 384] = 1'b1; frame0.error[ 384] = 1'b0;frame0.data[ 385] = 8'h74; frame0.valid[ 385] = 1'b1; frame0.error[ 385] = 1'b0;frame0.data[ 386] = 8'h75; frame0.valid[ 386] = 1'b1; frame0.error[ 386] = 1'b0;frame0.data[ 387] = 8'h76; frame0.valid[ 387] = 1'b1; frame0.error[ 387] = 1'b0;frame0.data[ 388] = 8'h77; frame0.valid[ 388] = 1'b1; frame0.error[ 388] = 1'b0;frame0.data[ 389] = 8'h78; frame0.valid[ 389] = 1'b1; frame0.error[ 389] = 1'b0;frame0.data[ 390] = 8'h79; frame0.valid[ 390] = 1'b1; frame0.error[ 390] = 1'b0;frame0.data[ 391] = 8'h7A; frame0.valid[ 391] = 1'b1; frame0.error[ 391] = 1'b0;frame0.data[ 392] = 8'h7B; frame0.valid[ 392] = 1'b1; frame0.error[ 392] = 1'b0;frame0.data[ 393] = 8'h7C; frame0.valid[ 393] = 1'b1; frame0.error[ 393] = 1'b0;frame0.data[ 394] = 8'h7D; frame0.valid[ 394] = 1'b1; frame0.error[ 394] = 1'b0;frame0.data[ 395] = 8'h7E; frame0.valid[ 395] = 1'b1; frame0.error[ 395] = 1'b0;frame0.data[ 396] = 8'h7F; frame0.valid[ 396] = 1'b1; frame0.error[ 396] = 1'b0;frame0.data[ 397] = 8'h80; frame0.valid[ 397] = 1'b1; frame0.error[ 397] = 1'b0;
        frame0.data[ 398] = 8'h81; frame0.valid[ 398] = 1'b1; frame0.error[ 398] = 1'b0;frame0.data[ 399] = 8'h82; frame0.valid[ 399] = 1'b1; frame0.error[ 399] = 1'b0;frame0.data[ 400] = 8'h83; frame0.valid[ 400] = 1'b1; frame0.error[ 400] = 1'b0;frame0.data[ 401] = 8'h84; frame0.valid[ 401] = 1'b1; frame0.error[ 401] = 1'b0;frame0.data[ 402] = 8'h85; frame0.valid[ 402] = 1'b1; frame0.error[ 402] = 1'b0;frame0.data[ 403] = 8'h86; frame0.valid[ 403] = 1'b1; frame0.error[ 403] = 1'b0;frame0.data[ 404] = 8'h87; frame0.valid[ 404] = 1'b1; frame0.error[ 404] = 1'b0;frame0.data[ 405] = 8'h88; frame0.valid[ 405] = 1'b1; frame0.error[ 405] = 1'b0;frame0.data[ 406] = 8'h89; frame0.valid[ 406] = 1'b1; frame0.error[ 406] = 1'b0;frame0.data[ 407] = 8'h8A; frame0.valid[ 407] = 1'b1; frame0.error[ 407] = 1'b0;frame0.data[ 408] = 8'h8B; frame0.valid[ 408] = 1'b1; frame0.error[ 408] = 1'b0;frame0.data[ 409] = 8'h8C; frame0.valid[ 409] = 1'b1; frame0.error[ 409] = 1'b0;frame0.data[ 410] = 8'h8D; frame0.valid[ 410] = 1'b1; frame0.error[ 410] = 1'b0;frame0.data[ 411] = 8'h8E; frame0.valid[ 411] = 1'b1; frame0.error[ 411] = 1'b0;frame0.data[ 412] = 8'h8F; frame0.valid[ 412] = 1'b1; frame0.error[ 412] = 1'b0;frame0.data[ 413] = 8'h90; frame0.valid[ 413] = 1'b1; frame0.error[ 413] = 1'b0;
        frame0.data[ 414] = 8'h91; frame0.valid[ 414] = 1'b1; frame0.error[ 414] = 1'b0;frame0.data[ 415] = 8'h92; frame0.valid[ 415] = 1'b1; frame0.error[ 415] = 1'b0;frame0.data[ 416] = 8'h93; frame0.valid[ 416] = 1'b1; frame0.error[ 416] = 1'b0;frame0.data[ 417] = 8'h94; frame0.valid[ 417] = 1'b1; frame0.error[ 417] = 1'b0;frame0.data[ 418] = 8'h95; frame0.valid[ 418] = 1'b1; frame0.error[ 418] = 1'b0;frame0.data[ 419] = 8'h96; frame0.valid[ 419] = 1'b1; frame0.error[ 419] = 1'b0;frame0.data[ 420] = 8'h97; frame0.valid[ 420] = 1'b1; frame0.error[ 420] = 1'b0;frame0.data[ 421] = 8'h98; frame0.valid[ 421] = 1'b1; frame0.error[ 421] = 1'b0;frame0.data[ 422] = 8'h99; frame0.valid[ 422] = 1'b1; frame0.error[ 422] = 1'b0;frame0.data[ 423] = 8'h9A; frame0.valid[ 423] = 1'b1; frame0.error[ 423] = 1'b0;frame0.data[ 424] = 8'h9B; frame0.valid[ 424] = 1'b1; frame0.error[ 424] = 1'b0;frame0.data[ 425] = 8'h9C; frame0.valid[ 425] = 1'b1; frame0.error[ 425] = 1'b0;frame0.data[ 426] = 8'h9D; frame0.valid[ 426] = 1'b1; frame0.error[ 426] = 1'b0;frame0.data[ 427] = 8'h9E; frame0.valid[ 427] = 1'b1; frame0.error[ 427] = 1'b0;frame0.data[ 428] = 8'h9F; frame0.valid[ 428] = 1'b1; frame0.error[ 428] = 1'b0;frame0.data[ 429] = 8'hA0; frame0.valid[ 429] = 1'b1; frame0.error[ 429] = 1'b0;
        frame0.data[ 430] = 8'hA1; frame0.valid[ 430] = 1'b1; frame0.error[ 430] = 1'b0;frame0.data[ 431] = 8'hA2; frame0.valid[ 431] = 1'b1; frame0.error[ 431] = 1'b0;frame0.data[ 432] = 8'hA3; frame0.valid[ 432] = 1'b1; frame0.error[ 432] = 1'b0;frame0.data[ 433] = 8'hA4; frame0.valid[ 433] = 1'b1; frame0.error[ 433] = 1'b0;frame0.data[ 434] = 8'hA5; frame0.valid[ 434] = 1'b1; frame0.error[ 434] = 1'b0;frame0.data[ 435] = 8'hA6; frame0.valid[ 435] = 1'b1; frame0.error[ 435] = 1'b0;frame0.data[ 436] = 8'hA7; frame0.valid[ 436] = 1'b1; frame0.error[ 436] = 1'b0;frame0.data[ 437] = 8'hA8; frame0.valid[ 437] = 1'b1; frame0.error[ 437] = 1'b0;frame0.data[ 438] = 8'hA9; frame0.valid[ 438] = 1'b1; frame0.error[ 438] = 1'b0;frame0.data[ 439] = 8'hAA; frame0.valid[ 439] = 1'b1; frame0.error[ 439] = 1'b0;frame0.data[ 440] = 8'hAB; frame0.valid[ 440] = 1'b1; frame0.error[ 440] = 1'b0;frame0.data[ 441] = 8'hAC; frame0.valid[ 441] = 1'b1; frame0.error[ 441] = 1'b0;frame0.data[ 442] = 8'hAD; frame0.valid[ 442] = 1'b1; frame0.error[ 442] = 1'b0;frame0.data[ 443] = 8'hAE; frame0.valid[ 443] = 1'b1; frame0.error[ 443] = 1'b0;frame0.data[ 444] = 8'hAF; frame0.valid[ 444] = 1'b1; frame0.error[ 444] = 1'b0;frame0.data[ 445] = 8'hB0; frame0.valid[ 445] = 1'b1; frame0.error[ 445] = 1'b0;
        frame0.data[ 446] = 8'hB1; frame0.valid[ 446] = 1'b1; frame0.error[ 446] = 1'b0;frame0.data[ 447] = 8'hB2; frame0.valid[ 447] = 1'b1; frame0.error[ 447] = 1'b0;frame0.data[ 448] = 8'hB3; frame0.valid[ 448] = 1'b1; frame0.error[ 448] = 1'b0;frame0.data[ 449] = 8'hB4; frame0.valid[ 449] = 1'b1; frame0.error[ 449] = 1'b0;frame0.data[ 450] = 8'hB5; frame0.valid[ 450] = 1'b1; frame0.error[ 450] = 1'b0;frame0.data[ 451] = 8'hB6; frame0.valid[ 451] = 1'b1; frame0.error[ 451] = 1'b0;frame0.data[ 452] = 8'hB7; frame0.valid[ 452] = 1'b1; frame0.error[ 452] = 1'b0;frame0.data[ 453] = 8'hB8; frame0.valid[ 453] = 1'b1; frame0.error[ 453] = 1'b0;frame0.data[ 454] = 8'hB9; frame0.valid[ 454] = 1'b1; frame0.error[ 454] = 1'b0;frame0.data[ 455] = 8'hBA; frame0.valid[ 455] = 1'b1; frame0.error[ 455] = 1'b0;frame0.data[ 456] = 8'hBB; frame0.valid[ 456] = 1'b1; frame0.error[ 456] = 1'b0;frame0.data[ 457] = 8'hBC; frame0.valid[ 457] = 1'b1; frame0.error[ 457] = 1'b0;frame0.data[ 458] = 8'hBD; frame0.valid[ 458] = 1'b1; frame0.error[ 458] = 1'b0;frame0.data[ 459] = 8'hBE; frame0.valid[ 459] = 1'b1; frame0.error[ 459] = 1'b0;frame0.data[ 460] = 8'hBF; frame0.valid[ 460] = 1'b1; frame0.error[ 460] = 1'b0;frame0.data[ 461] = 8'hC0; frame0.valid[ 461] = 1'b1; frame0.error[ 461] = 1'b0;
        frame0.data[ 462] = 8'hC1; frame0.valid[ 462] = 1'b1; frame0.error[ 462] = 1'b0;frame0.data[ 463] = 8'hC2; frame0.valid[ 463] = 1'b1; frame0.error[ 463] = 1'b0;frame0.data[ 464] = 8'hC3; frame0.valid[ 464] = 1'b1; frame0.error[ 464] = 1'b0;frame0.data[ 465] = 8'hC4; frame0.valid[ 465] = 1'b1; frame0.error[ 465] = 1'b0;frame0.data[ 466] = 8'hC5; frame0.valid[ 466] = 1'b1; frame0.error[ 466] = 1'b0;frame0.data[ 467] = 8'hC6; frame0.valid[ 467] = 1'b1; frame0.error[ 467] = 1'b0;frame0.data[ 468] = 8'hC7; frame0.valid[ 468] = 1'b1; frame0.error[ 468] = 1'b0;frame0.data[ 469] = 8'hC8; frame0.valid[ 469] = 1'b1; frame0.error[ 469] = 1'b0;frame0.data[ 470] = 8'hC9; frame0.valid[ 470] = 1'b1; frame0.error[ 470] = 1'b0;frame0.data[ 471] = 8'hCA; frame0.valid[ 471] = 1'b1; frame0.error[ 471] = 1'b0;frame0.data[ 472] = 8'hCB; frame0.valid[ 472] = 1'b1; frame0.error[ 472] = 1'b0;frame0.data[ 473] = 8'hCC; frame0.valid[ 473] = 1'b1; frame0.error[ 473] = 1'b0;frame0.data[ 474] = 8'hCD; frame0.valid[ 474] = 1'b1; frame0.error[ 474] = 1'b0;frame0.data[ 475] = 8'hCE; frame0.valid[ 475] = 1'b1; frame0.error[ 475] = 1'b0;frame0.data[ 476] = 8'hCF; frame0.valid[ 476] = 1'b1; frame0.error[ 476] = 1'b0;frame0.data[ 477] = 8'hD0; frame0.valid[ 477] = 1'b1; frame0.error[ 477] = 1'b0;
        frame0.data[ 478] = 8'hD1; frame0.valid[ 478] = 1'b1; frame0.error[ 478] = 1'b0;frame0.data[ 479] = 8'hD2; frame0.valid[ 479] = 1'b1; frame0.error[ 479] = 1'b0;frame0.data[ 480] = 8'hD3; frame0.valid[ 480] = 1'b1; frame0.error[ 480] = 1'b0;frame0.data[ 481] = 8'hD4; frame0.valid[ 481] = 1'b1; frame0.error[ 481] = 1'b0;frame0.data[ 482] = 8'hD5; frame0.valid[ 482] = 1'b1; frame0.error[ 482] = 1'b0;frame0.data[ 483] = 8'hD6; frame0.valid[ 483] = 1'b1; frame0.error[ 483] = 1'b0;frame0.data[ 484] = 8'hD7; frame0.valid[ 484] = 1'b1; frame0.error[ 484] = 1'b0;frame0.data[ 485] = 8'hD8; frame0.valid[ 485] = 1'b1; frame0.error[ 485] = 1'b0;frame0.data[ 486] = 8'hD9; frame0.valid[ 486] = 1'b1; frame0.error[ 486] = 1'b0;frame0.data[ 487] = 8'hDA; frame0.valid[ 487] = 1'b1; frame0.error[ 487] = 1'b0;frame0.data[ 488] = 8'hDB; frame0.valid[ 488] = 1'b1; frame0.error[ 488] = 1'b0;frame0.data[ 489] = 8'hDC; frame0.valid[ 489] = 1'b1; frame0.error[ 489] = 1'b0;frame0.data[ 490] = 8'hDD; frame0.valid[ 490] = 1'b1; frame0.error[ 490] = 1'b0;frame0.data[ 491] = 8'hDE; frame0.valid[ 491] = 1'b1; frame0.error[ 491] = 1'b0;frame0.data[ 492] = 8'hDF; frame0.valid[ 492] = 1'b1; frame0.error[ 492] = 1'b0;frame0.data[ 493] = 8'hE0; frame0.valid[ 493] = 1'b1; frame0.error[ 493] = 1'b0;
        frame0.data[ 494] = 8'hE1; frame0.valid[ 494] = 1'b1; frame0.error[ 494] = 1'b0;frame0.data[ 495] = 8'hE2; frame0.valid[ 495] = 1'b1; frame0.error[ 495] = 1'b0;frame0.data[ 496] = 8'hE3; frame0.valid[ 496] = 1'b1; frame0.error[ 496] = 1'b0;frame0.data[ 497] = 8'hE4; frame0.valid[ 497] = 1'b1; frame0.error[ 497] = 1'b0;frame0.data[ 498] = 8'hE5; frame0.valid[ 498] = 1'b1; frame0.error[ 498] = 1'b0;frame0.data[ 499] = 8'hE6; frame0.valid[ 499] = 1'b1; frame0.error[ 499] = 1'b0;frame0.data[ 500] = 8'hE7; frame0.valid[ 500] = 1'b1; frame0.error[ 500] = 1'b0;frame0.data[ 501] = 8'hE8; frame0.valid[ 501] = 1'b1; frame0.error[ 501] = 1'b0;frame0.data[ 502] = 8'hE9; frame0.valid[ 502] = 1'b1; frame0.error[ 502] = 1'b0;frame0.data[ 503] = 8'hEA; frame0.valid[ 503] = 1'b1; frame0.error[ 503] = 1'b0;frame0.data[ 504] = 8'hEB; frame0.valid[ 504] = 1'b1; frame0.error[ 504] = 1'b0;frame0.data[ 505] = 8'hEC; frame0.valid[ 505] = 1'b1; frame0.error[ 505] = 1'b0;frame0.data[ 506] = 8'hED; frame0.valid[ 506] = 1'b1; frame0.error[ 506] = 1'b0;frame0.data[ 507] = 8'hEE; frame0.valid[ 507] = 1'b1; frame0.error[ 507] = 1'b0;frame0.data[ 508] = 8'hEF; frame0.valid[ 508] = 1'b1; frame0.error[ 508] = 1'b0;frame0.data[ 509] = 8'hF0; frame0.valid[ 509] = 1'b1; frame0.error[ 509] = 1'b0;
        frame0.data[ 510] = 8'hF1; frame0.valid[ 510] = 1'b1; frame0.error[ 510] = 1'b0;frame0.data[ 511] = 8'hF2; frame0.valid[ 511] = 1'b1; frame0.error[ 511] = 1'b0;frame0.data[ 512] = 8'hF3; frame0.valid[ 512] = 1'b1; frame0.error[ 512] = 1'b0;frame0.data[ 513] = 8'hF4; frame0.valid[ 513] = 1'b1; frame0.error[ 513] = 1'b0;frame0.data[ 514] = 8'hF5; frame0.valid[ 514] = 1'b1; frame0.error[ 514] = 1'b0;frame0.data[ 515] = 8'hF6; frame0.valid[ 515] = 1'b1; frame0.error[ 515] = 1'b0;frame0.data[ 516] = 8'hF7; frame0.valid[ 516] = 1'b1; frame0.error[ 516] = 1'b0;frame0.data[ 517] = 8'hF8; frame0.valid[ 517] = 1'b1; frame0.error[ 517] = 1'b0;frame0.data[ 518] = 8'hF9; frame0.valid[ 518] = 1'b1; frame0.error[ 518] = 1'b0;frame0.data[ 519] = 8'hFA; frame0.valid[ 519] = 1'b1; frame0.error[ 519] = 1'b0;frame0.data[ 520] = 8'hFB; frame0.valid[ 520] = 1'b1; frame0.error[ 520] = 1'b0;frame0.data[ 521] = 8'hFC; frame0.valid[ 521] = 1'b1; frame0.error[ 521] = 1'b0;frame0.data[ 522] = 8'hFD; frame0.valid[ 522] = 1'b1; frame0.error[ 522] = 1'b0;frame0.data[ 523] = 8'hFE; frame0.valid[ 523] = 1'b1; frame0.error[ 523] = 1'b0;frame0.data[ 524] = 8'h00; frame0.valid[ 524] = 1'b1; frame0.error[ 524] = 1'b0;frame0.data[ 525] = 8'h01; frame0.valid[ 525] = 1'b1; frame0.error[ 525] = 1'b0;
        frame0.data[ 526] = 8'h02; frame0.valid[ 526] = 1'b1; frame0.error[ 526] = 1'b0;frame0.data[ 527] = 8'h03; frame0.valid[ 527] = 1'b1; frame0.error[ 527] = 1'b0;frame0.data[ 528] = 8'h04; frame0.valid[ 528] = 1'b1; frame0.error[ 528] = 1'b0;frame0.data[ 529] = 8'h05; frame0.valid[ 529] = 1'b1; frame0.error[ 529] = 1'b0;frame0.data[ 530] = 8'h06; frame0.valid[ 530] = 1'b1; frame0.error[ 530] = 1'b0;frame0.data[ 531] = 8'h07; frame0.valid[ 531] = 1'b1; frame0.error[ 531] = 1'b0;frame0.data[ 532] = 8'h08; frame0.valid[ 532] = 1'b1; frame0.error[ 532] = 1'b0;frame0.data[ 533] = 8'h09; frame0.valid[ 533] = 1'b1; frame0.error[ 533] = 1'b0;frame0.data[ 534] = 8'h0A; frame0.valid[ 534] = 1'b1; frame0.error[ 534] = 1'b0;frame0.data[ 535] = 8'h0B; frame0.valid[ 535] = 1'b1; frame0.error[ 535] = 1'b0;frame0.data[ 536] = 8'h0C; frame0.valid[ 536] = 1'b1; frame0.error[ 536] = 1'b0;frame0.data[ 537] = 8'h0D; frame0.valid[ 537] = 1'b1; frame0.error[ 537] = 1'b0;frame0.data[ 538] = 8'h0E; frame0.valid[ 538] = 1'b1; frame0.error[ 538] = 1'b0;frame0.data[ 539] = 8'h0F; frame0.valid[ 539] = 1'b1; frame0.error[ 539] = 1'b0;frame0.data[ 540] = 8'h10; frame0.valid[ 540] = 1'b1; frame0.error[ 540] = 1'b0;frame0.data[ 541] = 8'h11; frame0.valid[ 541] = 1'b1; frame0.error[ 541] = 1'b0;
        frame0.data[ 542] = 8'h12; frame0.valid[ 542] = 1'b1; frame0.error[ 542] = 1'b0;frame0.data[ 543] = 8'h13; frame0.valid[ 543] = 1'b1; frame0.error[ 543] = 1'b0;frame0.data[ 544] = 8'h14; frame0.valid[ 544] = 1'b1; frame0.error[ 544] = 1'b0;frame0.data[ 545] = 8'h15; frame0.valid[ 545] = 1'b1; frame0.error[ 545] = 1'b0;frame0.data[ 546] = 8'h16; frame0.valid[ 546] = 1'b1; frame0.error[ 546] = 1'b0;frame0.data[ 547] = 8'h17; frame0.valid[ 547] = 1'b1; frame0.error[ 547] = 1'b0;frame0.data[ 548] = 8'h18; frame0.valid[ 548] = 1'b1; frame0.error[ 548] = 1'b0;frame0.data[ 549] = 8'h19; frame0.valid[ 549] = 1'b1; frame0.error[ 549] = 1'b0;frame0.data[ 550] = 8'h1A; frame0.valid[ 550] = 1'b1; frame0.error[ 550] = 1'b0;frame0.data[ 551] = 8'h1B; frame0.valid[ 551] = 1'b1; frame0.error[ 551] = 1'b0;frame0.data[ 552] = 8'h1C; frame0.valid[ 552] = 1'b1; frame0.error[ 552] = 1'b0;frame0.data[ 553] = 8'h1D; frame0.valid[ 553] = 1'b1; frame0.error[ 553] = 1'b0;frame0.data[ 554] = 8'h1E; frame0.valid[ 554] = 1'b1; frame0.error[ 554] = 1'b0;frame0.data[ 555] = 8'h1F; frame0.valid[ 555] = 1'b1; frame0.error[ 555] = 1'b0;frame0.data[ 556] = 8'h20; frame0.valid[ 556] = 1'b1; frame0.error[ 556] = 1'b0;frame0.data[ 557] = 8'h21; frame0.valid[ 557] = 1'b1; frame0.error[ 557] = 1'b0;
        frame0.data[ 558] = 8'h22; frame0.valid[ 558] = 1'b1; frame0.error[ 558] = 1'b0;frame0.data[ 559] = 8'h23; frame0.valid[ 559] = 1'b1; frame0.error[ 559] = 1'b0;frame0.data[ 560] = 8'h24; frame0.valid[ 560] = 1'b1; frame0.error[ 560] = 1'b0;frame0.data[ 561] = 8'h25; frame0.valid[ 561] = 1'b1; frame0.error[ 561] = 1'b0;frame0.data[ 562] = 8'h26; frame0.valid[ 562] = 1'b1; frame0.error[ 562] = 1'b0;frame0.data[ 563] = 8'h27; frame0.valid[ 563] = 1'b1; frame0.error[ 563] = 1'b0;frame0.data[ 564] = 8'h28; frame0.valid[ 564] = 1'b1; frame0.error[ 564] = 1'b0;frame0.data[ 565] = 8'h29; frame0.valid[ 565] = 1'b1; frame0.error[ 565] = 1'b0;frame0.data[ 566] = 8'h2A; frame0.valid[ 566] = 1'b1; frame0.error[ 566] = 1'b0;frame0.data[ 567] = 8'h2B; frame0.valid[ 567] = 1'b1; frame0.error[ 567] = 1'b0;frame0.data[ 568] = 8'h2C; frame0.valid[ 568] = 1'b1; frame0.error[ 568] = 1'b0;frame0.data[ 569] = 8'h2D; frame0.valid[ 569] = 1'b1; frame0.error[ 569] = 1'b0;frame0.data[ 570] = 8'h2E; frame0.valid[ 570] = 1'b1; frame0.error[ 570] = 1'b0;frame0.data[ 571] = 8'h2F; frame0.valid[ 571] = 1'b1; frame0.error[ 571] = 1'b0;frame0.data[ 572] = 8'h30; frame0.valid[ 572] = 1'b1; frame0.error[ 572] = 1'b0;frame0.data[ 573] = 8'h31; frame0.valid[ 573] = 1'b1; frame0.error[ 573] = 1'b0;
        frame0.data[ 574] = 8'h32; frame0.valid[ 574] = 1'b1; frame0.error[ 574] = 1'b0;frame0.data[ 575] = 8'h33; frame0.valid[ 575] = 1'b1; frame0.error[ 575] = 1'b0;frame0.data[ 576] = 8'h34; frame0.valid[ 576] = 1'b1; frame0.error[ 576] = 1'b0;frame0.data[ 577] = 8'h35; frame0.valid[ 577] = 1'b1; frame0.error[ 577] = 1'b0;frame0.data[ 578] = 8'h36; frame0.valid[ 578] = 1'b1; frame0.error[ 578] = 1'b0;frame0.data[ 579] = 8'h37; frame0.valid[ 579] = 1'b1; frame0.error[ 579] = 1'b0;frame0.data[ 580] = 8'h38; frame0.valid[ 580] = 1'b1; frame0.error[ 580] = 1'b0;frame0.data[ 581] = 8'h39; frame0.valid[ 581] = 1'b1; frame0.error[ 581] = 1'b0;frame0.data[ 582] = 8'h3A; frame0.valid[ 582] = 1'b1; frame0.error[ 582] = 1'b0;frame0.data[ 583] = 8'h3B; frame0.valid[ 583] = 1'b1; frame0.error[ 583] = 1'b0;frame0.data[ 584] = 8'h3C; frame0.valid[ 584] = 1'b1; frame0.error[ 584] = 1'b0;frame0.data[ 585] = 8'h3D; frame0.valid[ 585] = 1'b1; frame0.error[ 585] = 1'b0;frame0.data[ 586] = 8'h3E; frame0.valid[ 586] = 1'b1; frame0.error[ 586] = 1'b0;frame0.data[ 587] = 8'h3F; frame0.valid[ 587] = 1'b1; frame0.error[ 587] = 1'b0;frame0.data[ 588] = 8'h40; frame0.valid[ 588] = 1'b1; frame0.error[ 588] = 1'b0;frame0.data[ 589] = 8'h41; frame0.valid[ 589] = 1'b1; frame0.error[ 589] = 1'b0;
        frame0.data[ 590] = 8'h42; frame0.valid[ 590] = 1'b1; frame0.error[ 590] = 1'b0;frame0.data[ 591] = 8'h43; frame0.valid[ 591] = 1'b1; frame0.error[ 591] = 1'b0;frame0.data[ 592] = 8'h44; frame0.valid[ 592] = 1'b1; frame0.error[ 592] = 1'b0;frame0.data[ 593] = 8'h45; frame0.valid[ 593] = 1'b1; frame0.error[ 593] = 1'b0;frame0.data[ 594] = 8'h46; frame0.valid[ 594] = 1'b1; frame0.error[ 594] = 1'b0;frame0.data[ 595] = 8'h47; frame0.valid[ 595] = 1'b1; frame0.error[ 595] = 1'b0;frame0.data[ 596] = 8'h48; frame0.valid[ 596] = 1'b1; frame0.error[ 596] = 1'b0;frame0.data[ 597] = 8'h49; frame0.valid[ 597] = 1'b1; frame0.error[ 597] = 1'b0;frame0.data[ 598] = 8'h4A; frame0.valid[ 598] = 1'b1; frame0.error[ 598] = 1'b0;frame0.data[ 599] = 8'h4B; frame0.valid[ 599] = 1'b1; frame0.error[ 599] = 1'b0;frame0.data[ 600] = 8'h4C; frame0.valid[ 600] = 1'b1; frame0.error[ 600] = 1'b0;frame0.data[ 601] = 8'h4D; frame0.valid[ 601] = 1'b1; frame0.error[ 601] = 1'b0;frame0.data[ 602] = 8'h4E; frame0.valid[ 602] = 1'b1; frame0.error[ 602] = 1'b0;frame0.data[ 603] = 8'h4F; frame0.valid[ 603] = 1'b1; frame0.error[ 603] = 1'b0;frame0.data[ 604] = 8'h50; frame0.valid[ 604] = 1'b1; frame0.error[ 604] = 1'b0;frame0.data[ 605] = 8'h51; frame0.valid[ 605] = 1'b1; frame0.error[ 605] = 1'b0;
        frame0.data[ 606] = 8'h52; frame0.valid[ 606] = 1'b1; frame0.error[ 606] = 1'b0;frame0.data[ 607] = 8'h53; frame0.valid[ 607] = 1'b1; frame0.error[ 607] = 1'b0;frame0.data[ 608] = 8'h54; frame0.valid[ 608] = 1'b1; frame0.error[ 608] = 1'b0;frame0.data[ 609] = 8'h55; frame0.valid[ 609] = 1'b1; frame0.error[ 609] = 1'b0;frame0.data[ 610] = 8'h56; frame0.valid[ 610] = 1'b1; frame0.error[ 610] = 1'b0;frame0.data[ 611] = 8'h57; frame0.valid[ 611] = 1'b1; frame0.error[ 611] = 1'b0;frame0.data[ 612] = 8'h58; frame0.valid[ 612] = 1'b1; frame0.error[ 612] = 1'b0;frame0.data[ 613] = 8'h59; frame0.valid[ 613] = 1'b1; frame0.error[ 613] = 1'b0;frame0.data[ 614] = 8'h5A; frame0.valid[ 614] = 1'b1; frame0.error[ 614] = 1'b0;frame0.data[ 615] = 8'h5B; frame0.valid[ 615] = 1'b1; frame0.error[ 615] = 1'b0;frame0.data[ 616] = 8'h5C; frame0.valid[ 616] = 1'b1; frame0.error[ 616] = 1'b0;frame0.data[ 617] = 8'h5D; frame0.valid[ 617] = 1'b1; frame0.error[ 617] = 1'b0;frame0.data[ 618] = 8'h5E; frame0.valid[ 618] = 1'b1; frame0.error[ 618] = 1'b0;frame0.data[ 619] = 8'h5F; frame0.valid[ 619] = 1'b1; frame0.error[ 619] = 1'b0;frame0.data[ 620] = 8'h60; frame0.valid[ 620] = 1'b1; frame0.error[ 620] = 1'b0;frame0.data[ 621] = 8'h61; frame0.valid[ 621] = 1'b1; frame0.error[ 621] = 1'b0;
        frame0.data[ 622] = 8'h62; frame0.valid[ 622] = 1'b1; frame0.error[ 622] = 1'b0;frame0.data[ 623] = 8'h63; frame0.valid[ 623] = 1'b1; frame0.error[ 623] = 1'b0;frame0.data[ 624] = 8'h64; frame0.valid[ 624] = 1'b1; frame0.error[ 624] = 1'b0;frame0.data[ 625] = 8'h65; frame0.valid[ 625] = 1'b1; frame0.error[ 625] = 1'b0;frame0.data[ 626] = 8'h66; frame0.valid[ 626] = 1'b1; frame0.error[ 626] = 1'b0;frame0.data[ 627] = 8'h67; frame0.valid[ 627] = 1'b1; frame0.error[ 627] = 1'b0;frame0.data[ 628] = 8'h68; frame0.valid[ 628] = 1'b1; frame0.error[ 628] = 1'b0;frame0.data[ 629] = 8'h69; frame0.valid[ 629] = 1'b1; frame0.error[ 629] = 1'b0;frame0.data[ 630] = 8'h6A; frame0.valid[ 630] = 1'b1; frame0.error[ 630] = 1'b0;frame0.data[ 631] = 8'h6B; frame0.valid[ 631] = 1'b1; frame0.error[ 631] = 1'b0;frame0.data[ 632] = 8'h6C; frame0.valid[ 632] = 1'b1; frame0.error[ 632] = 1'b0;frame0.data[ 633] = 8'h6D; frame0.valid[ 633] = 1'b1; frame0.error[ 633] = 1'b0;frame0.data[ 634] = 8'h6E; frame0.valid[ 634] = 1'b1; frame0.error[ 634] = 1'b0;frame0.data[ 635] = 8'h6F; frame0.valid[ 635] = 1'b1; frame0.error[ 635] = 1'b0;frame0.data[ 636] = 8'h70; frame0.valid[ 636] = 1'b1; frame0.error[ 636] = 1'b0;frame0.data[ 637] = 8'h71; frame0.valid[ 637] = 1'b1; frame0.error[ 637] = 1'b0;
        frame0.data[ 638] = 8'h72; frame0.valid[ 638] = 1'b1; frame0.error[ 638] = 1'b0;frame0.data[ 639] = 8'h73; frame0.valid[ 639] = 1'b1; frame0.error[ 639] = 1'b0;frame0.data[ 640] = 8'h74; frame0.valid[ 640] = 1'b1; frame0.error[ 640] = 1'b0;frame0.data[ 641] = 8'h75; frame0.valid[ 641] = 1'b1; frame0.error[ 641] = 1'b0;frame0.data[ 642] = 8'h76; frame0.valid[ 642] = 1'b1; frame0.error[ 642] = 1'b0;frame0.data[ 643] = 8'h77; frame0.valid[ 643] = 1'b1; frame0.error[ 643] = 1'b0;frame0.data[ 644] = 8'h78; frame0.valid[ 644] = 1'b1; frame0.error[ 644] = 1'b0;frame0.data[ 645] = 8'h79; frame0.valid[ 645] = 1'b1; frame0.error[ 645] = 1'b0;frame0.data[ 646] = 8'h7A; frame0.valid[ 646] = 1'b1; frame0.error[ 646] = 1'b0;frame0.data[ 647] = 8'h7B; frame0.valid[ 647] = 1'b1; frame0.error[ 647] = 1'b0;frame0.data[ 648] = 8'h7C; frame0.valid[ 648] = 1'b1; frame0.error[ 648] = 1'b0;frame0.data[ 649] = 8'h7D; frame0.valid[ 649] = 1'b1; frame0.error[ 649] = 1'b0;frame0.data[ 650] = 8'h7E; frame0.valid[ 650] = 1'b1; frame0.error[ 650] = 1'b0;frame0.data[ 651] = 8'h7F; frame0.valid[ 651] = 1'b1; frame0.error[ 651] = 1'b0;frame0.data[ 652] = 8'h80; frame0.valid[ 652] = 1'b1; frame0.error[ 652] = 1'b0;frame0.data[ 653] = 8'h81; frame0.valid[ 653] = 1'b1; frame0.error[ 653] = 1'b0;
        frame0.data[ 654] = 8'h82; frame0.valid[ 654] = 1'b1; frame0.error[ 654] = 1'b0;frame0.data[ 655] = 8'h83; frame0.valid[ 655] = 1'b1; frame0.error[ 655] = 1'b0;frame0.data[ 656] = 8'h84; frame0.valid[ 656] = 1'b1; frame0.error[ 656] = 1'b0;frame0.data[ 657] = 8'h85; frame0.valid[ 657] = 1'b1; frame0.error[ 657] = 1'b0;frame0.data[ 658] = 8'h86; frame0.valid[ 658] = 1'b1; frame0.error[ 658] = 1'b0;frame0.data[ 659] = 8'h87; frame0.valid[ 659] = 1'b1; frame0.error[ 659] = 1'b0;frame0.data[ 660] = 8'h88; frame0.valid[ 660] = 1'b1; frame0.error[ 660] = 1'b0;frame0.data[ 661] = 8'h89; frame0.valid[ 661] = 1'b1; frame0.error[ 661] = 1'b0;frame0.data[ 662] = 8'h8A; frame0.valid[ 662] = 1'b1; frame0.error[ 662] = 1'b0;frame0.data[ 663] = 8'h8B; frame0.valid[ 663] = 1'b1; frame0.error[ 663] = 1'b0;frame0.data[ 664] = 8'h8C; frame0.valid[ 664] = 1'b1; frame0.error[ 664] = 1'b0;frame0.data[ 665] = 8'h8D; frame0.valid[ 665] = 1'b1; frame0.error[ 665] = 1'b0;frame0.data[ 666] = 8'h8E; frame0.valid[ 666] = 1'b1; frame0.error[ 666] = 1'b0;frame0.data[ 667] = 8'h8F; frame0.valid[ 667] = 1'b1; frame0.error[ 667] = 1'b0;frame0.data[ 668] = 8'h90; frame0.valid[ 668] = 1'b1; frame0.error[ 668] = 1'b0;frame0.data[ 669] = 8'h91; frame0.valid[ 669] = 1'b1; frame0.error[ 669] = 1'b0;
        frame0.data[ 670] = 8'h92; frame0.valid[ 670] = 1'b1; frame0.error[ 670] = 1'b0;frame0.data[ 671] = 8'h93; frame0.valid[ 671] = 1'b1; frame0.error[ 671] = 1'b0;frame0.data[ 672] = 8'h94; frame0.valid[ 672] = 1'b1; frame0.error[ 672] = 1'b0;frame0.data[ 673] = 8'h95; frame0.valid[ 673] = 1'b1; frame0.error[ 673] = 1'b0;frame0.data[ 674] = 8'h96; frame0.valid[ 674] = 1'b1; frame0.error[ 674] = 1'b0;frame0.data[ 675] = 8'h97; frame0.valid[ 675] = 1'b1; frame0.error[ 675] = 1'b0;frame0.data[ 676] = 8'h98; frame0.valid[ 676] = 1'b1; frame0.error[ 676] = 1'b0;frame0.data[ 677] = 8'h99; frame0.valid[ 677] = 1'b1; frame0.error[ 677] = 1'b0;frame0.data[ 678] = 8'h9A; frame0.valid[ 678] = 1'b1; frame0.error[ 678] = 1'b0;frame0.data[ 679] = 8'h9B; frame0.valid[ 679] = 1'b1; frame0.error[ 679] = 1'b0;frame0.data[ 680] = 8'h9C; frame0.valid[ 680] = 1'b1; frame0.error[ 680] = 1'b0;frame0.data[ 681] = 8'h9D; frame0.valid[ 681] = 1'b1; frame0.error[ 681] = 1'b0;frame0.data[ 682] = 8'h9E; frame0.valid[ 682] = 1'b1; frame0.error[ 682] = 1'b0;frame0.data[ 683] = 8'h9F; frame0.valid[ 683] = 1'b1; frame0.error[ 683] = 1'b0;frame0.data[ 684] = 8'hA0; frame0.valid[ 684] = 1'b1; frame0.error[ 684] = 1'b0;frame0.data[ 685] = 8'hA1; frame0.valid[ 685] = 1'b1; frame0.error[ 685] = 1'b0;
        frame0.data[ 686] = 8'hA2; frame0.valid[ 686] = 1'b1; frame0.error[ 686] = 1'b0;frame0.data[ 687] = 8'hA3; frame0.valid[ 687] = 1'b1; frame0.error[ 687] = 1'b0;frame0.data[ 688] = 8'hA4; frame0.valid[ 688] = 1'b1; frame0.error[ 688] = 1'b0;frame0.data[ 689] = 8'hA5; frame0.valid[ 689] = 1'b1; frame0.error[ 689] = 1'b0;frame0.data[ 690] = 8'hA6; frame0.valid[ 690] = 1'b1; frame0.error[ 690] = 1'b0;frame0.data[ 691] = 8'hA7; frame0.valid[ 691] = 1'b1; frame0.error[ 691] = 1'b0;frame0.data[ 692] = 8'hA8; frame0.valid[ 692] = 1'b1; frame0.error[ 692] = 1'b0;frame0.data[ 693] = 8'hA9; frame0.valid[ 693] = 1'b1; frame0.error[ 693] = 1'b0;frame0.data[ 694] = 8'hAA; frame0.valid[ 694] = 1'b1; frame0.error[ 694] = 1'b0;frame0.data[ 695] = 8'hAB; frame0.valid[ 695] = 1'b1; frame0.error[ 695] = 1'b0;frame0.data[ 696] = 8'hAC; frame0.valid[ 696] = 1'b1; frame0.error[ 696] = 1'b0;frame0.data[ 697] = 8'hAD; frame0.valid[ 697] = 1'b1; frame0.error[ 697] = 1'b0;frame0.data[ 698] = 8'hAE; frame0.valid[ 698] = 1'b1; frame0.error[ 698] = 1'b0;frame0.data[ 699] = 8'hAF; frame0.valid[ 699] = 1'b1; frame0.error[ 699] = 1'b0;frame0.data[ 700] = 8'hB0; frame0.valid[ 700] = 1'b1; frame0.error[ 700] = 1'b0;frame0.data[ 701] = 8'hB1; frame0.valid[ 701] = 1'b1; frame0.error[ 701] = 1'b0;
        frame0.data[ 702] = 8'hB2; frame0.valid[ 702] = 1'b1; frame0.error[ 702] = 1'b0;frame0.data[ 703] = 8'hB3; frame0.valid[ 703] = 1'b1; frame0.error[ 703] = 1'b0;frame0.data[ 704] = 8'hB4; frame0.valid[ 704] = 1'b1; frame0.error[ 704] = 1'b0;frame0.data[ 705] = 8'hB5; frame0.valid[ 705] = 1'b1; frame0.error[ 705] = 1'b0;frame0.data[ 706] = 8'hB6; frame0.valid[ 706] = 1'b1; frame0.error[ 706] = 1'b0;frame0.data[ 707] = 8'hB7; frame0.valid[ 707] = 1'b1; frame0.error[ 707] = 1'b0;frame0.data[ 708] = 8'hB8; frame0.valid[ 708] = 1'b1; frame0.error[ 708] = 1'b0;frame0.data[ 709] = 8'hB9; frame0.valid[ 709] = 1'b1; frame0.error[ 709] = 1'b0;frame0.data[ 710] = 8'hBA; frame0.valid[ 710] = 1'b1; frame0.error[ 710] = 1'b0;frame0.data[ 711] = 8'hBB; frame0.valid[ 711] = 1'b1; frame0.error[ 711] = 1'b0;frame0.data[ 712] = 8'hBC; frame0.valid[ 712] = 1'b1; frame0.error[ 712] = 1'b0;frame0.data[ 713] = 8'hBD; frame0.valid[ 713] = 1'b1; frame0.error[ 713] = 1'b0;frame0.data[ 714] = 8'hBE; frame0.valid[ 714] = 1'b1; frame0.error[ 714] = 1'b0;frame0.data[ 715] = 8'hBF; frame0.valid[ 715] = 1'b1; frame0.error[ 715] = 1'b0;frame0.data[ 716] = 8'hC0; frame0.valid[ 716] = 1'b1; frame0.error[ 716] = 1'b0;frame0.data[ 717] = 8'hC1; frame0.valid[ 717] = 1'b1; frame0.error[ 717] = 1'b0;
        frame0.data[ 718] = 8'hC2; frame0.valid[ 718] = 1'b1; frame0.error[ 718] = 1'b0;frame0.data[ 719] = 8'hC3; frame0.valid[ 719] = 1'b1; frame0.error[ 719] = 1'b0;frame0.data[ 720] = 8'hC4; frame0.valid[ 720] = 1'b1; frame0.error[ 720] = 1'b0;frame0.data[ 721] = 8'hC5; frame0.valid[ 721] = 1'b1; frame0.error[ 721] = 1'b0;frame0.data[ 722] = 8'hC6; frame0.valid[ 722] = 1'b1; frame0.error[ 722] = 1'b0;frame0.data[ 723] = 8'hC7; frame0.valid[ 723] = 1'b1; frame0.error[ 723] = 1'b0;frame0.data[ 724] = 8'hC8; frame0.valid[ 724] = 1'b1; frame0.error[ 724] = 1'b0;frame0.data[ 725] = 8'hC9; frame0.valid[ 725] = 1'b1; frame0.error[ 725] = 1'b0;frame0.data[ 726] = 8'hCA; frame0.valid[ 726] = 1'b1; frame0.error[ 726] = 1'b0;frame0.data[ 727] = 8'hCB; frame0.valid[ 727] = 1'b1; frame0.error[ 727] = 1'b0;frame0.data[ 728] = 8'hCC; frame0.valid[ 728] = 1'b1; frame0.error[ 728] = 1'b0;frame0.data[ 729] = 8'hCD; frame0.valid[ 729] = 1'b1; frame0.error[ 729] = 1'b0;frame0.data[ 730] = 8'hCE; frame0.valid[ 730] = 1'b1; frame0.error[ 730] = 1'b0;frame0.data[ 731] = 8'hCF; frame0.valid[ 731] = 1'b1; frame0.error[ 731] = 1'b0;frame0.data[ 732] = 8'hD0; frame0.valid[ 732] = 1'b1; frame0.error[ 732] = 1'b0;frame0.data[ 733] = 8'hD1; frame0.valid[ 733] = 1'b1; frame0.error[ 733] = 1'b0;
        frame0.data[ 734] = 8'hD2; frame0.valid[ 734] = 1'b1; frame0.error[ 734] = 1'b0;frame0.data[ 735] = 8'hD3; frame0.valid[ 735] = 1'b1; frame0.error[ 735] = 1'b0;frame0.data[ 736] = 8'hD4; frame0.valid[ 736] = 1'b1; frame0.error[ 736] = 1'b0;frame0.data[ 737] = 8'hD5; frame0.valid[ 737] = 1'b1; frame0.error[ 737] = 1'b0;frame0.data[ 738] = 8'hD6; frame0.valid[ 738] = 1'b1; frame0.error[ 738] = 1'b0;frame0.data[ 739] = 8'hD7; frame0.valid[ 739] = 1'b1; frame0.error[ 739] = 1'b0;frame0.data[ 740] = 8'hD8; frame0.valid[ 740] = 1'b1; frame0.error[ 740] = 1'b0;frame0.data[ 741] = 8'hD9; frame0.valid[ 741] = 1'b1; frame0.error[ 741] = 1'b0;frame0.data[ 742] = 8'hDA; frame0.valid[ 742] = 1'b1; frame0.error[ 742] = 1'b0;frame0.data[ 743] = 8'hDB; frame0.valid[ 743] = 1'b1; frame0.error[ 743] = 1'b0;frame0.data[ 744] = 8'hDC; frame0.valid[ 744] = 1'b1; frame0.error[ 744] = 1'b0;frame0.data[ 745] = 8'hDD; frame0.valid[ 745] = 1'b1; frame0.error[ 745] = 1'b0;frame0.data[ 746] = 8'hDE; frame0.valid[ 746] = 1'b1; frame0.error[ 746] = 1'b0;frame0.data[ 747] = 8'hDF; frame0.valid[ 747] = 1'b1; frame0.error[ 747] = 1'b0;frame0.data[ 748] = 8'hE0; frame0.valid[ 748] = 1'b1; frame0.error[ 748] = 1'b0;frame0.data[ 749] = 8'hE1; frame0.valid[ 749] = 1'b1; frame0.error[ 749] = 1'b0;
        frame0.data[ 750] = 8'hE2; frame0.valid[ 750] = 1'b1; frame0.error[ 750] = 1'b0;frame0.data[ 751] = 8'hE3; frame0.valid[ 751] = 1'b1; frame0.error[ 751] = 1'b0;frame0.data[ 752] = 8'hE4; frame0.valid[ 752] = 1'b1; frame0.error[ 752] = 1'b0;frame0.data[ 753] = 8'hE5; frame0.valid[ 753] = 1'b1; frame0.error[ 753] = 1'b0;frame0.data[ 754] = 8'hE6; frame0.valid[ 754] = 1'b1; frame0.error[ 754] = 1'b0;frame0.data[ 755] = 8'hE7; frame0.valid[ 755] = 1'b1; frame0.error[ 755] = 1'b0;frame0.data[ 756] = 8'hE8; frame0.valid[ 756] = 1'b1; frame0.error[ 756] = 1'b0;frame0.data[ 757] = 8'hE9; frame0.valid[ 757] = 1'b1; frame0.error[ 757] = 1'b0;frame0.data[ 758] = 8'hEA; frame0.valid[ 758] = 1'b1; frame0.error[ 758] = 1'b0;frame0.data[ 759] = 8'hEB; frame0.valid[ 759] = 1'b1; frame0.error[ 759] = 1'b0;frame0.data[ 760] = 8'hEC; frame0.valid[ 760] = 1'b1; frame0.error[ 760] = 1'b0;frame0.data[ 761] = 8'hED; frame0.valid[ 761] = 1'b1; frame0.error[ 761] = 1'b0;frame0.data[ 762] = 8'hEE; frame0.valid[ 762] = 1'b1; frame0.error[ 762] = 1'b0;frame0.data[ 763] = 8'hEF; frame0.valid[ 763] = 1'b1; frame0.error[ 763] = 1'b0;frame0.data[ 764] = 8'hF0; frame0.valid[ 764] = 1'b1; frame0.error[ 764] = 1'b0;frame0.data[ 765] = 8'hF1; frame0.valid[ 765] = 1'b1; frame0.error[ 765] = 1'b0;
        frame0.data[ 766] = 8'hF2; frame0.valid[ 766] = 1'b1; frame0.error[ 766] = 1'b0;frame0.data[ 767] = 8'hF3; frame0.valid[ 767] = 1'b1; frame0.error[ 767] = 1'b0;frame0.data[ 768] = 8'hF4; frame0.valid[ 768] = 1'b1; frame0.error[ 768] = 1'b0;frame0.data[ 769] = 8'hF5; frame0.valid[ 769] = 1'b1; frame0.error[ 769] = 1'b0;frame0.data[ 770] = 8'hF6; frame0.valid[ 770] = 1'b1; frame0.error[ 770] = 1'b0;frame0.data[ 771] = 8'hF7; frame0.valid[ 771] = 1'b1; frame0.error[ 771] = 1'b0;frame0.data[ 772] = 8'hF8; frame0.valid[ 772] = 1'b1; frame0.error[ 772] = 1'b0;frame0.data[ 773] = 8'hF9; frame0.valid[ 773] = 1'b1; frame0.error[ 773] = 1'b0;frame0.data[ 774] = 8'hFA; frame0.valid[ 774] = 1'b1; frame0.error[ 774] = 1'b0;frame0.data[ 775] = 8'hFB; frame0.valid[ 775] = 1'b1; frame0.error[ 775] = 1'b0;frame0.data[ 776] = 8'hFC; frame0.valid[ 776] = 1'b1; frame0.error[ 776] = 1'b0;frame0.data[ 777] = 8'hFD; frame0.valid[ 777] = 1'b1; frame0.error[ 777] = 1'b0;frame0.data[ 778] = 8'hFE; frame0.valid[ 778] = 1'b1; frame0.error[ 778] = 1'b0;frame0.data[ 779] = 8'h00; frame0.valid[ 779] = 1'b1; frame0.error[ 779] = 1'b0;frame0.data[ 780] = 8'h01; frame0.valid[ 780] = 1'b1; frame0.error[ 780] = 1'b0;frame0.data[ 781] = 8'h02; frame0.valid[ 781] = 1'b1; frame0.error[ 781] = 1'b0;
        frame0.data[ 782] = 8'h03; frame0.valid[ 782] = 1'b1; frame0.error[ 782] = 1'b0;frame0.data[ 783] = 8'h04; frame0.valid[ 783] = 1'b1; frame0.error[ 783] = 1'b0;frame0.data[ 784] = 8'h05; frame0.valid[ 784] = 1'b1; frame0.error[ 784] = 1'b0;frame0.data[ 785] = 8'h06; frame0.valid[ 785] = 1'b1; frame0.error[ 785] = 1'b0;frame0.data[ 786] = 8'h07; frame0.valid[ 786] = 1'b1; frame0.error[ 786] = 1'b0;frame0.data[ 787] = 8'h08; frame0.valid[ 787] = 1'b1; frame0.error[ 787] = 1'b0;frame0.data[ 788] = 8'h09; frame0.valid[ 788] = 1'b1; frame0.error[ 788] = 1'b0;frame0.data[ 789] = 8'h0A; frame0.valid[ 789] = 1'b1; frame0.error[ 789] = 1'b0;frame0.data[ 790] = 8'h0B; frame0.valid[ 790] = 1'b1; frame0.error[ 790] = 1'b0;frame0.data[ 791] = 8'h0C; frame0.valid[ 791] = 1'b1; frame0.error[ 791] = 1'b0;frame0.data[ 792] = 8'h0D; frame0.valid[ 792] = 1'b1; frame0.error[ 792] = 1'b0;frame0.data[ 793] = 8'h0E; frame0.valid[ 793] = 1'b1; frame0.error[ 793] = 1'b0;frame0.data[ 794] = 8'h0F; frame0.valid[ 794] = 1'b1; frame0.error[ 794] = 1'b0;frame0.data[ 795] = 8'h10; frame0.valid[ 795] = 1'b1; frame0.error[ 795] = 1'b0;frame0.data[ 796] = 8'h11; frame0.valid[ 796] = 1'b1; frame0.error[ 796] = 1'b0;frame0.data[ 797] = 8'h12; frame0.valid[ 797] = 1'b1; frame0.error[ 797] = 1'b0;
        frame0.data[ 798] = 8'h13; frame0.valid[ 798] = 1'b1; frame0.error[ 798] = 1'b0;frame0.data[ 799] = 8'h14; frame0.valid[ 799] = 1'b1; frame0.error[ 799] = 1'b0;frame0.data[ 800] = 8'h15; frame0.valid[ 800] = 1'b1; frame0.error[ 800] = 1'b0;frame0.data[ 801] = 8'h16; frame0.valid[ 801] = 1'b1; frame0.error[ 801] = 1'b0;frame0.data[ 802] = 8'h17; frame0.valid[ 802] = 1'b1; frame0.error[ 802] = 1'b0;frame0.data[ 803] = 8'h18; frame0.valid[ 803] = 1'b1; frame0.error[ 803] = 1'b0;frame0.data[ 804] = 8'h19; frame0.valid[ 804] = 1'b1; frame0.error[ 804] = 1'b0;frame0.data[ 805] = 8'h1A; frame0.valid[ 805] = 1'b1; frame0.error[ 805] = 1'b0;frame0.data[ 806] = 8'h1B; frame0.valid[ 806] = 1'b1; frame0.error[ 806] = 1'b0;frame0.data[ 807] = 8'h1C; frame0.valid[ 807] = 1'b1; frame0.error[ 807] = 1'b0;frame0.data[ 808] = 8'h1D; frame0.valid[ 808] = 1'b1; frame0.error[ 808] = 1'b0;frame0.data[ 809] = 8'h1E; frame0.valid[ 809] = 1'b1; frame0.error[ 809] = 1'b0;frame0.data[ 810] = 8'h1F; frame0.valid[ 810] = 1'b1; frame0.error[ 810] = 1'b0;frame0.data[ 811] = 8'h20; frame0.valid[ 811] = 1'b1; frame0.error[ 811] = 1'b0;frame0.data[ 812] = 8'h21; frame0.valid[ 812] = 1'b1; frame0.error[ 812] = 1'b0;frame0.data[ 813] = 8'h22; frame0.valid[ 813] = 1'b1; frame0.error[ 813] = 1'b0;
        frame0.data[ 814] = 8'h23; frame0.valid[ 814] = 1'b1; frame0.error[ 814] = 1'b0;frame0.data[ 815] = 8'h24; frame0.valid[ 815] = 1'b1; frame0.error[ 815] = 1'b0;frame0.data[ 816] = 8'h25; frame0.valid[ 816] = 1'b1; frame0.error[ 816] = 1'b0;frame0.data[ 817] = 8'h26; frame0.valid[ 817] = 1'b1; frame0.error[ 817] = 1'b0;frame0.data[ 818] = 8'h27; frame0.valid[ 818] = 1'b1; frame0.error[ 818] = 1'b0;frame0.data[ 819] = 8'h28; frame0.valid[ 819] = 1'b1; frame0.error[ 819] = 1'b0;frame0.data[ 820] = 8'h29; frame0.valid[ 820] = 1'b1; frame0.error[ 820] = 1'b0;frame0.data[ 821] = 8'h2A; frame0.valid[ 821] = 1'b1; frame0.error[ 821] = 1'b0;frame0.data[ 822] = 8'h2B; frame0.valid[ 822] = 1'b1; frame0.error[ 822] = 1'b0;frame0.data[ 823] = 8'h2C; frame0.valid[ 823] = 1'b1; frame0.error[ 823] = 1'b0;frame0.data[ 824] = 8'h2D; frame0.valid[ 824] = 1'b1; frame0.error[ 824] = 1'b0;frame0.data[ 825] = 8'h2E; frame0.valid[ 825] = 1'b1; frame0.error[ 825] = 1'b0;frame0.data[ 826] = 8'h2F; frame0.valid[ 826] = 1'b1; frame0.error[ 826] = 1'b0;frame0.data[ 827] = 8'h30; frame0.valid[ 827] = 1'b1; frame0.error[ 827] = 1'b0;frame0.data[ 828] = 8'h31; frame0.valid[ 828] = 1'b1; frame0.error[ 828] = 1'b0;frame0.data[ 829] = 8'h32; frame0.valid[ 829] = 1'b1; frame0.error[ 829] = 1'b0;
        frame0.data[ 830] = 8'h33; frame0.valid[ 830] = 1'b1; frame0.error[ 830] = 1'b0;frame0.data[ 831] = 8'h34; frame0.valid[ 831] = 1'b1; frame0.error[ 831] = 1'b0;frame0.data[ 832] = 8'h35; frame0.valid[ 832] = 1'b1; frame0.error[ 832] = 1'b0;frame0.data[ 833] = 8'h36; frame0.valid[ 833] = 1'b1; frame0.error[ 833] = 1'b0;frame0.data[ 834] = 8'h37; frame0.valid[ 834] = 1'b1; frame0.error[ 834] = 1'b0;frame0.data[ 835] = 8'h38; frame0.valid[ 835] = 1'b1; frame0.error[ 835] = 1'b0;frame0.data[ 836] = 8'h39; frame0.valid[ 836] = 1'b1; frame0.error[ 836] = 1'b0;frame0.data[ 837] = 8'h3A; frame0.valid[ 837] = 1'b1; frame0.error[ 837] = 1'b0;frame0.data[ 838] = 8'h3B; frame0.valid[ 838] = 1'b1; frame0.error[ 838] = 1'b0;frame0.data[ 839] = 8'h3C; frame0.valid[ 839] = 1'b1; frame0.error[ 839] = 1'b0;frame0.data[ 840] = 8'h3D; frame0.valid[ 840] = 1'b1; frame0.error[ 840] = 1'b0;frame0.data[ 841] = 8'h3E; frame0.valid[ 841] = 1'b1; frame0.error[ 841] = 1'b0;frame0.data[ 842] = 8'h3F; frame0.valid[ 842] = 1'b1; frame0.error[ 842] = 1'b0;frame0.data[ 843] = 8'h40; frame0.valid[ 843] = 1'b1; frame0.error[ 843] = 1'b0;frame0.data[ 844] = 8'h41; frame0.valid[ 844] = 1'b1; frame0.error[ 844] = 1'b0;frame0.data[ 845] = 8'h42; frame0.valid[ 845] = 1'b1; frame0.error[ 845] = 1'b0;
        frame0.data[ 846] = 8'h43; frame0.valid[ 846] = 1'b1; frame0.error[ 846] = 1'b0;frame0.data[ 847] = 8'h44; frame0.valid[ 847] = 1'b1; frame0.error[ 847] = 1'b0;frame0.data[ 848] = 8'h45; frame0.valid[ 848] = 1'b1; frame0.error[ 848] = 1'b0;frame0.data[ 849] = 8'h46; frame0.valid[ 849] = 1'b1; frame0.error[ 849] = 1'b0;frame0.data[ 850] = 8'h47; frame0.valid[ 850] = 1'b1; frame0.error[ 850] = 1'b0;frame0.data[ 851] = 8'h48; frame0.valid[ 851] = 1'b1; frame0.error[ 851] = 1'b0;frame0.data[ 852] = 8'h49; frame0.valid[ 852] = 1'b1; frame0.error[ 852] = 1'b0;frame0.data[ 853] = 8'h4A; frame0.valid[ 853] = 1'b1; frame0.error[ 853] = 1'b0;frame0.data[ 854] = 8'h4B; frame0.valid[ 854] = 1'b1; frame0.error[ 854] = 1'b0;frame0.data[ 855] = 8'h4C; frame0.valid[ 855] = 1'b1; frame0.error[ 855] = 1'b0;frame0.data[ 856] = 8'h4D; frame0.valid[ 856] = 1'b1; frame0.error[ 856] = 1'b0;frame0.data[ 857] = 8'h4E; frame0.valid[ 857] = 1'b1; frame0.error[ 857] = 1'b0;frame0.data[ 858] = 8'h4F; frame0.valid[ 858] = 1'b1; frame0.error[ 858] = 1'b0;frame0.data[ 859] = 8'h50; frame0.valid[ 859] = 1'b1; frame0.error[ 859] = 1'b0;frame0.data[ 860] = 8'h51; frame0.valid[ 860] = 1'b1; frame0.error[ 860] = 1'b0;frame0.data[ 861] = 8'h52; frame0.valid[ 861] = 1'b1; frame0.error[ 861] = 1'b0;
        frame0.data[ 862] = 8'h53; frame0.valid[ 862] = 1'b1; frame0.error[ 862] = 1'b0;frame0.data[ 863] = 8'h54; frame0.valid[ 863] = 1'b1; frame0.error[ 863] = 1'b0;frame0.data[ 864] = 8'h55; frame0.valid[ 864] = 1'b1; frame0.error[ 864] = 1'b0;frame0.data[ 865] = 8'h56; frame0.valid[ 865] = 1'b1; frame0.error[ 865] = 1'b0;frame0.data[ 866] = 8'h57; frame0.valid[ 866] = 1'b1; frame0.error[ 866] = 1'b0;frame0.data[ 867] = 8'h58; frame0.valid[ 867] = 1'b1; frame0.error[ 867] = 1'b0;frame0.data[ 868] = 8'h59; frame0.valid[ 868] = 1'b1; frame0.error[ 868] = 1'b0;frame0.data[ 869] = 8'h5A; frame0.valid[ 869] = 1'b1; frame0.error[ 869] = 1'b0;frame0.data[ 870] = 8'h5B; frame0.valid[ 870] = 1'b1; frame0.error[ 870] = 1'b0;frame0.data[ 871] = 8'h5C; frame0.valid[ 871] = 1'b1; frame0.error[ 871] = 1'b0;frame0.data[ 872] = 8'h5D; frame0.valid[ 872] = 1'b1; frame0.error[ 872] = 1'b0;frame0.data[ 873] = 8'h5E; frame0.valid[ 873] = 1'b1; frame0.error[ 873] = 1'b0;frame0.data[ 874] = 8'h5F; frame0.valid[ 874] = 1'b1; frame0.error[ 874] = 1'b0;frame0.data[ 875] = 8'h60; frame0.valid[ 875] = 1'b1; frame0.error[ 875] = 1'b0;frame0.data[ 876] = 8'h61; frame0.valid[ 876] = 1'b1; frame0.error[ 876] = 1'b0;frame0.data[ 877] = 8'h62; frame0.valid[ 877] = 1'b1; frame0.error[ 877] = 1'b0;
        frame0.data[ 878] = 8'h63; frame0.valid[ 878] = 1'b1; frame0.error[ 878] = 1'b0;frame0.data[ 879] = 8'h64; frame0.valid[ 879] = 1'b1; frame0.error[ 879] = 1'b0;frame0.data[ 880] = 8'h65; frame0.valid[ 880] = 1'b1; frame0.error[ 880] = 1'b0;frame0.data[ 881] = 8'h66; frame0.valid[ 881] = 1'b1; frame0.error[ 881] = 1'b0;frame0.data[ 882] = 8'h67; frame0.valid[ 882] = 1'b1; frame0.error[ 882] = 1'b0;frame0.data[ 883] = 8'h68; frame0.valid[ 883] = 1'b1; frame0.error[ 883] = 1'b0;frame0.data[ 884] = 8'h69; frame0.valid[ 884] = 1'b1; frame0.error[ 884] = 1'b0;frame0.data[ 885] = 8'h6A; frame0.valid[ 885] = 1'b1; frame0.error[ 885] = 1'b0;frame0.data[ 886] = 8'h6B; frame0.valid[ 886] = 1'b1; frame0.error[ 886] = 1'b0;frame0.data[ 887] = 8'h6C; frame0.valid[ 887] = 1'b1; frame0.error[ 887] = 1'b0;frame0.data[ 888] = 8'h6D; frame0.valid[ 888] = 1'b1; frame0.error[ 888] = 1'b0;frame0.data[ 889] = 8'h6E; frame0.valid[ 889] = 1'b1; frame0.error[ 889] = 1'b0;frame0.data[ 890] = 8'h6F; frame0.valid[ 890] = 1'b1; frame0.error[ 890] = 1'b0;frame0.data[ 891] = 8'h70; frame0.valid[ 891] = 1'b1; frame0.error[ 891] = 1'b0;frame0.data[ 892] = 8'h71; frame0.valid[ 892] = 1'b1; frame0.error[ 892] = 1'b0;frame0.data[ 893] = 8'h72; frame0.valid[ 893] = 1'b1; frame0.error[ 893] = 1'b0;
        frame0.data[ 894] = 8'h73; frame0.valid[ 894] = 1'b1; frame0.error[ 894] = 1'b0;frame0.data[ 895] = 8'h74; frame0.valid[ 895] = 1'b1; frame0.error[ 895] = 1'b0;frame0.data[ 896] = 8'h75; frame0.valid[ 896] = 1'b1; frame0.error[ 896] = 1'b0;frame0.data[ 897] = 8'h76; frame0.valid[ 897] = 1'b1; frame0.error[ 897] = 1'b0;frame0.data[ 898] = 8'h77; frame0.valid[ 898] = 1'b1; frame0.error[ 898] = 1'b0;frame0.data[ 899] = 8'h78; frame0.valid[ 899] = 1'b1; frame0.error[ 899] = 1'b0;frame0.data[ 900] = 8'h79; frame0.valid[ 900] = 1'b1; frame0.error[ 900] = 1'b0;frame0.data[ 901] = 8'h7A; frame0.valid[ 901] = 1'b1; frame0.error[ 901] = 1'b0;frame0.data[ 902] = 8'h7B; frame0.valid[ 902] = 1'b1; frame0.error[ 902] = 1'b0;frame0.data[ 903] = 8'h7C; frame0.valid[ 903] = 1'b1; frame0.error[ 903] = 1'b0;frame0.data[ 904] = 8'h7D; frame0.valid[ 904] = 1'b1; frame0.error[ 904] = 1'b0;frame0.data[ 905] = 8'h7E; frame0.valid[ 905] = 1'b1; frame0.error[ 905] = 1'b0;frame0.data[ 906] = 8'h7F; frame0.valid[ 906] = 1'b1; frame0.error[ 906] = 1'b0;frame0.data[ 907] = 8'h80; frame0.valid[ 907] = 1'b1; frame0.error[ 907] = 1'b0;frame0.data[ 908] = 8'h81; frame0.valid[ 908] = 1'b1; frame0.error[ 908] = 1'b0;frame0.data[ 909] = 8'h82; frame0.valid[ 909] = 1'b1; frame0.error[ 909] = 1'b0;
        frame0.data[ 910] = 8'h83; frame0.valid[ 910] = 1'b1; frame0.error[ 910] = 1'b0;frame0.data[ 911] = 8'h84; frame0.valid[ 911] = 1'b1; frame0.error[ 911] = 1'b0;frame0.data[ 912] = 8'h85; frame0.valid[ 912] = 1'b1; frame0.error[ 912] = 1'b0;frame0.data[ 913] = 8'h86; frame0.valid[ 913] = 1'b1; frame0.error[ 913] = 1'b0;frame0.data[ 914] = 8'h87; frame0.valid[ 914] = 1'b1; frame0.error[ 914] = 1'b0;frame0.data[ 915] = 8'h88; frame0.valid[ 915] = 1'b1; frame0.error[ 915] = 1'b0;frame0.data[ 916] = 8'h89; frame0.valid[ 916] = 1'b1; frame0.error[ 916] = 1'b0;frame0.data[ 917] = 8'h8A; frame0.valid[ 917] = 1'b1; frame0.error[ 917] = 1'b0;frame0.data[ 918] = 8'h8B; frame0.valid[ 918] = 1'b1; frame0.error[ 918] = 1'b0;frame0.data[ 919] = 8'h8C; frame0.valid[ 919] = 1'b1; frame0.error[ 919] = 1'b0;frame0.data[ 920] = 8'h8D; frame0.valid[ 920] = 1'b1; frame0.error[ 920] = 1'b0;frame0.data[ 921] = 8'h8E; frame0.valid[ 921] = 1'b1; frame0.error[ 921] = 1'b0;frame0.data[ 922] = 8'h8F; frame0.valid[ 922] = 1'b1; frame0.error[ 922] = 1'b0;frame0.data[ 923] = 8'h90; frame0.valid[ 923] = 1'b1; frame0.error[ 923] = 1'b0;frame0.data[ 924] = 8'h91; frame0.valid[ 924] = 1'b1; frame0.error[ 924] = 1'b0;frame0.data[ 925] = 8'h92; frame0.valid[ 925] = 1'b1; frame0.error[ 925] = 1'b0;
        frame0.data[ 926] = 8'h93; frame0.valid[ 926] = 1'b1; frame0.error[ 926] = 1'b0;frame0.data[ 927] = 8'h94; frame0.valid[ 927] = 1'b1; frame0.error[ 927] = 1'b0;frame0.data[ 928] = 8'h95; frame0.valid[ 928] = 1'b1; frame0.error[ 928] = 1'b0;frame0.data[ 929] = 8'h96; frame0.valid[ 929] = 1'b1; frame0.error[ 929] = 1'b0;frame0.data[ 930] = 8'h97; frame0.valid[ 930] = 1'b1; frame0.error[ 930] = 1'b0;frame0.data[ 931] = 8'h98; frame0.valid[ 931] = 1'b1; frame0.error[ 931] = 1'b0;frame0.data[ 932] = 8'h99; frame0.valid[ 932] = 1'b1; frame0.error[ 932] = 1'b0;frame0.data[ 933] = 8'h9A; frame0.valid[ 933] = 1'b1; frame0.error[ 933] = 1'b0;frame0.data[ 934] = 8'h9B; frame0.valid[ 934] = 1'b1; frame0.error[ 934] = 1'b0;frame0.data[ 935] = 8'h9C; frame0.valid[ 935] = 1'b1; frame0.error[ 935] = 1'b0;frame0.data[ 936] = 8'h9D; frame0.valid[ 936] = 1'b1; frame0.error[ 936] = 1'b0;frame0.data[ 937] = 8'h9E; frame0.valid[ 937] = 1'b1; frame0.error[ 937] = 1'b0;frame0.data[ 938] = 8'h9F; frame0.valid[ 938] = 1'b1; frame0.error[ 938] = 1'b0;frame0.data[ 939] = 8'hA0; frame0.valid[ 939] = 1'b1; frame0.error[ 939] = 1'b0;frame0.data[ 940] = 8'hA1; frame0.valid[ 940] = 1'b1; frame0.error[ 940] = 1'b0;frame0.data[ 941] = 8'hA2; frame0.valid[ 941] = 1'b1; frame0.error[ 941] = 1'b0;
        frame0.data[ 942] = 8'hA3; frame0.valid[ 942] = 1'b1; frame0.error[ 942] = 1'b0;frame0.data[ 943] = 8'hA4; frame0.valid[ 943] = 1'b1; frame0.error[ 943] = 1'b0;frame0.data[ 944] = 8'hA5; frame0.valid[ 944] = 1'b1; frame0.error[ 944] = 1'b0;frame0.data[ 945] = 8'hA6; frame0.valid[ 945] = 1'b1; frame0.error[ 945] = 1'b0;frame0.data[ 946] = 8'hA7; frame0.valid[ 946] = 1'b1; frame0.error[ 946] = 1'b0;frame0.data[ 947] = 8'hA8; frame0.valid[ 947] = 1'b1; frame0.error[ 947] = 1'b0;frame0.data[ 948] = 8'hA9; frame0.valid[ 948] = 1'b1; frame0.error[ 948] = 1'b0;frame0.data[ 949] = 8'hAA; frame0.valid[ 949] = 1'b1; frame0.error[ 949] = 1'b0;frame0.data[ 950] = 8'hAB; frame0.valid[ 950] = 1'b1; frame0.error[ 950] = 1'b0;frame0.data[ 951] = 8'hAC; frame0.valid[ 951] = 1'b1; frame0.error[ 951] = 1'b0;frame0.data[ 952] = 8'hAD; frame0.valid[ 952] = 1'b1; frame0.error[ 952] = 1'b0;frame0.data[ 953] = 8'hAE; frame0.valid[ 953] = 1'b1; frame0.error[ 953] = 1'b0;frame0.data[ 954] = 8'hAF; frame0.valid[ 954] = 1'b1; frame0.error[ 954] = 1'b0;frame0.data[ 955] = 8'hB0; frame0.valid[ 955] = 1'b1; frame0.error[ 955] = 1'b0;frame0.data[ 956] = 8'hB1; frame0.valid[ 956] = 1'b1; frame0.error[ 956] = 1'b0;frame0.data[ 957] = 8'hB2; frame0.valid[ 957] = 1'b1; frame0.error[ 957] = 1'b0;
        frame0.data[ 958] = 8'hB3; frame0.valid[ 958] = 1'b1; frame0.error[ 958] = 1'b0;frame0.data[ 959] = 8'hB4; frame0.valid[ 959] = 1'b1; frame0.error[ 959] = 1'b0;frame0.data[ 960] = 8'hB5; frame0.valid[ 960] = 1'b1; frame0.error[ 960] = 1'b0;frame0.data[ 961] = 8'hB6; frame0.valid[ 961] = 1'b1; frame0.error[ 961] = 1'b0;frame0.data[ 962] = 8'hB7; frame0.valid[ 962] = 1'b1; frame0.error[ 962] = 1'b0;frame0.data[ 963] = 8'hB8; frame0.valid[ 963] = 1'b1; frame0.error[ 963] = 1'b0;frame0.data[ 964] = 8'hB9; frame0.valid[ 964] = 1'b1; frame0.error[ 964] = 1'b0;frame0.data[ 965] = 8'hBA; frame0.valid[ 965] = 1'b1; frame0.error[ 965] = 1'b0;frame0.data[ 966] = 8'hBB; frame0.valid[ 966] = 1'b1; frame0.error[ 966] = 1'b0;frame0.data[ 967] = 8'hBC; frame0.valid[ 967] = 1'b1; frame0.error[ 967] = 1'b0;frame0.data[ 968] = 8'hBD; frame0.valid[ 968] = 1'b1; frame0.error[ 968] = 1'b0;frame0.data[ 969] = 8'hBE; frame0.valid[ 969] = 1'b1; frame0.error[ 969] = 1'b0;frame0.data[ 970] = 8'hBF; frame0.valid[ 970] = 1'b1; frame0.error[ 970] = 1'b0;frame0.data[ 971] = 8'hC0; frame0.valid[ 971] = 1'b1; frame0.error[ 971] = 1'b0;frame0.data[ 972] = 8'hC1; frame0.valid[ 972] = 1'b1; frame0.error[ 972] = 1'b0;frame0.data[ 973] = 8'hC2; frame0.valid[ 973] = 1'b1; frame0.error[ 973] = 1'b0;
        frame0.data[ 974] = 8'hC3; frame0.valid[ 974] = 1'b1; frame0.error[ 974] = 1'b0;frame0.data[ 975] = 8'hC4; frame0.valid[ 975] = 1'b1; frame0.error[ 975] = 1'b0;frame0.data[ 976] = 8'hC5; frame0.valid[ 976] = 1'b1; frame0.error[ 976] = 1'b0;frame0.data[ 977] = 8'hC6; frame0.valid[ 977] = 1'b1; frame0.error[ 977] = 1'b0;frame0.data[ 978] = 8'hC7; frame0.valid[ 978] = 1'b1; frame0.error[ 978] = 1'b0;frame0.data[ 979] = 8'hC8; frame0.valid[ 979] = 1'b1; frame0.error[ 979] = 1'b0;frame0.data[ 980] = 8'hC9; frame0.valid[ 980] = 1'b1; frame0.error[ 980] = 1'b0;frame0.data[ 981] = 8'hCA; frame0.valid[ 981] = 1'b1; frame0.error[ 981] = 1'b0;frame0.data[ 982] = 8'hCB; frame0.valid[ 982] = 1'b1; frame0.error[ 982] = 1'b0;frame0.data[ 983] = 8'hCC; frame0.valid[ 983] = 1'b1; frame0.error[ 983] = 1'b0;frame0.data[ 984] = 8'hCD; frame0.valid[ 984] = 1'b1; frame0.error[ 984] = 1'b0;frame0.data[ 985] = 8'hCE; frame0.valid[ 985] = 1'b1; frame0.error[ 985] = 1'b0;frame0.data[ 986] = 8'hCF; frame0.valid[ 986] = 1'b1; frame0.error[ 986] = 1'b0;frame0.data[ 987] = 8'hD0; frame0.valid[ 987] = 1'b1; frame0.error[ 987] = 1'b0;frame0.data[ 988] = 8'hD1; frame0.valid[ 988] = 1'b1; frame0.error[ 988] = 1'b0;frame0.data[ 989] = 8'hD2; frame0.valid[ 989] = 1'b1; frame0.error[ 989] = 1'b0;
        frame0.data[ 990] = 8'hD3; frame0.valid[ 990] = 1'b1; frame0.error[ 990] = 1'b0;frame0.data[ 991] = 8'hD4; frame0.valid[ 991] = 1'b1; frame0.error[ 991] = 1'b0;frame0.data[ 992] = 8'hD5; frame0.valid[ 992] = 1'b1; frame0.error[ 992] = 1'b0;frame0.data[ 993] = 8'hD6; frame0.valid[ 993] = 1'b1; frame0.error[ 993] = 1'b0;frame0.data[ 994] = 8'hD7; frame0.valid[ 994] = 1'b1; frame0.error[ 994] = 1'b0;frame0.data[ 995] = 8'hD8; frame0.valid[ 995] = 1'b1; frame0.error[ 995] = 1'b0;frame0.data[ 996] = 8'hD9; frame0.valid[ 996] = 1'b1; frame0.error[ 996] = 1'b0;frame0.data[ 997] = 8'hDA; frame0.valid[ 997] = 1'b1; frame0.error[ 997] = 1'b0;frame0.data[ 998] = 8'hDB; frame0.valid[ 998] = 1'b1; frame0.error[ 998] = 1'b0;frame0.data[ 999] = 8'hDC; frame0.valid[ 999] = 1'b1; frame0.error[ 999] = 1'b0;frame0.data[1000] = 8'hDD; frame0.valid[1000] = 1'b1; frame0.error[1000] = 1'b0;frame0.data[1001] = 8'hDE; frame0.valid[1001] = 1'b1; frame0.error[1001] = 1'b0;frame0.data[1002] = 8'hDF; frame0.valid[1002] = 1'b1; frame0.error[1002] = 1'b0;frame0.data[1003] = 8'hE0; frame0.valid[1003] = 1'b1; frame0.error[1003] = 1'b0;frame0.data[1004] = 8'hE1; frame0.valid[1004] = 1'b1; frame0.error[1004] = 1'b0;frame0.data[1005] = 8'hE2; frame0.valid[1005] = 1'b1; frame0.error[1005] = 1'b0;
        frame0.data[1006] = 8'hE3; frame0.valid[1006] = 1'b1; frame0.error[1006] = 1'b0;frame0.data[1007] = 8'hE4; frame0.valid[1007] = 1'b1; frame0.error[1007] = 1'b0;frame0.data[1008] = 8'hE5; frame0.valid[1008] = 1'b1; frame0.error[1008] = 1'b0;frame0.data[1009] = 8'hE6; frame0.valid[1009] = 1'b1; frame0.error[1009] = 1'b0;frame0.data[1010] = 8'hE7; frame0.valid[1010] = 1'b1; frame0.error[1010] = 1'b0;frame0.data[1011] = 8'hE8; frame0.valid[1011] = 1'b1; frame0.error[1011] = 1'b0;frame0.data[1012] = 8'hE9; frame0.valid[1012] = 1'b1; frame0.error[1012] = 1'b0;frame0.data[1013] = 8'hEA; frame0.valid[1013] = 1'b1; frame0.error[1013] = 1'b0;frame0.data[1014] = 8'hEB; frame0.valid[1014] = 1'b1; frame0.error[1014] = 1'b0;frame0.data[1015] = 8'hEC; frame0.valid[1015] = 1'b1; frame0.error[1015] = 1'b0;frame0.data[1016] = 8'hED; frame0.valid[1016] = 1'b1; frame0.error[1016] = 1'b0;frame0.data[1017] = 8'hEE; frame0.valid[1017] = 1'b1; frame0.error[1017] = 1'b0;frame0.data[1018] = 8'hEF; frame0.valid[1018] = 1'b1; frame0.error[1018] = 1'b0;frame0.data[1019] = 8'hF0; frame0.valid[1019] = 1'b1; frame0.error[1019] = 1'b0;frame0.data[1020] = 8'hF1; frame0.valid[1020] = 1'b1; frame0.error[1020] = 1'b0;frame0.data[1021] = 8'hF2; frame0.valid[1021] = 1'b1; frame0.error[1021] = 1'b0;
        frame0.data[1022] = 8'hF3; frame0.valid[1022] = 1'b1; frame0.error[1022] = 1'b0;frame0.data[1023] = 8'hF4; frame0.valid[1023] = 1'b1; frame0.error[1023] = 1'b0;frame0.data[1024] = 8'hF5; frame0.valid[1024] = 1'b1; frame0.error[1024] = 1'b0;frame0.data[1025] = 8'hF6; frame0.valid[1025] = 1'b1; frame0.error[1025] = 1'b0;frame0.data[1026] = 8'hF7; frame0.valid[1026] = 1'b1; frame0.error[1026] = 1'b0;frame0.data[1027] = 8'hF8; frame0.valid[1027] = 1'b1; frame0.error[1027] = 1'b0;frame0.data[1028] = 8'hF9; frame0.valid[1028] = 1'b1; frame0.error[1028] = 1'b0;frame0.data[1029] = 8'hFA; frame0.valid[1029] = 1'b1; frame0.error[1029] = 1'b0;frame0.data[1030] = 8'hFB; frame0.valid[1030] = 1'b1; frame0.error[1030] = 1'b0;frame0.data[1031] = 8'hFC; frame0.valid[1031] = 1'b1; frame0.error[1031] = 1'b0;frame0.data[1032] = 8'hFD; frame0.valid[1032] = 1'b1; frame0.error[1032] = 1'b0;frame0.data[1033] = 8'hFE; frame0.valid[1033] = 1'b1; frame0.error[1033] = 1'b0;frame0.data[1034] = 8'h00; frame0.valid[1034] = 1'b1; frame0.error[1034] = 1'b0;frame0.data[1035] = 8'h01; frame0.valid[1035] = 1'b1; frame0.error[1035] = 1'b0;frame0.data[1036] = 8'h02; frame0.valid[1036] = 1'b1; frame0.error[1036] = 1'b0;frame0.data[1037] = 8'h03; frame0.valid[1037] = 1'b1; frame0.error[1037] = 1'b0;
        frame0.data[1038] = 8'h04; frame0.valid[1038] = 1'b1; frame0.error[1038] = 1'b0;frame0.data[1039] = 8'h05; frame0.valid[1039] = 1'b1; frame0.error[1039] = 1'b0;frame0.data[1040] = 8'h06; frame0.valid[1040] = 1'b1; frame0.error[1040] = 1'b0;frame0.data[1041] = 8'h07; frame0.valid[1041] = 1'b1; frame0.error[1041] = 1'b0;frame0.data[1042] = 8'h08; frame0.valid[1042] = 1'b1; frame0.error[1042] = 1'b0;frame0.data[1043] = 8'h09; frame0.valid[1043] = 1'b1; frame0.error[1043] = 1'b0;frame0.data[1044] = 8'h0A; frame0.valid[1044] = 1'b1; frame0.error[1044] = 1'b0;frame0.data[1045] = 8'h0B; frame0.valid[1045] = 1'b1; frame0.error[1045] = 1'b0;frame0.data[1046] = 8'h0C; frame0.valid[1046] = 1'b1; frame0.error[1046] = 1'b0;frame0.data[1047] = 8'h0D; frame0.valid[1047] = 1'b1; frame0.error[1047] = 1'b0;frame0.data[1048] = 8'h0E; frame0.valid[1048] = 1'b1; frame0.error[1048] = 1'b0;frame0.data[1049] = 8'h0F; frame0.valid[1049] = 1'b1; frame0.error[1049] = 1'b0;frame0.data[1050] = 8'h10; frame0.valid[1050] = 1'b1; frame0.error[1050] = 1'b0;frame0.data[1051] = 8'h11; frame0.valid[1051] = 1'b1; frame0.error[1051] = 1'b0;frame0.data[1052] = 8'h12; frame0.valid[1052] = 1'b1; frame0.error[1052] = 1'b0;frame0.data[1053] = 8'h13; frame0.valid[1053] = 1'b1; frame0.error[1053] = 1'b0;
        frame0.data[1054] = 8'h14; frame0.valid[1054] = 1'b1; frame0.error[1054] = 1'b0;frame0.data[1055] = 8'h15; frame0.valid[1055] = 1'b1; frame0.error[1055] = 1'b0;frame0.data[1056] = 8'h16; frame0.valid[1056] = 1'b1; frame0.error[1056] = 1'b0;frame0.data[1057] = 8'h17; frame0.valid[1057] = 1'b1; frame0.error[1057] = 1'b0;frame0.data[1058] = 8'h18; frame0.valid[1058] = 1'b1; frame0.error[1058] = 1'b0;frame0.data[1059] = 8'h19; frame0.valid[1059] = 1'b1; frame0.error[1059] = 1'b0;frame0.data[1060] = 8'h1A; frame0.valid[1060] = 1'b1; frame0.error[1060] = 1'b0;frame0.data[1061] = 8'h1B; frame0.valid[1061] = 1'b1; frame0.error[1061] = 1'b0;frame0.data[1062] = 8'h1C; frame0.valid[1062] = 1'b1; frame0.error[1062] = 1'b0;frame0.data[1063] = 8'h1D; frame0.valid[1063] = 1'b1; frame0.error[1063] = 1'b0;frame0.data[1064] = 8'h1E; frame0.valid[1064] = 1'b1; frame0.error[1064] = 1'b0;frame0.data[1065] = 8'h1F; frame0.valid[1065] = 1'b1; frame0.error[1065] = 1'b0;frame0.data[1066] = 8'h20; frame0.valid[1066] = 1'b1; frame0.error[1066] = 1'b0;frame0.data[1067] = 8'h21; frame0.valid[1067] = 1'b1; frame0.error[1067] = 1'b0;frame0.data[1068] = 8'h22; frame0.valid[1068] = 1'b1; frame0.error[1068] = 1'b0;frame0.data[1069] = 8'h23; frame0.valid[1069] = 1'b1; frame0.error[1069] = 1'b0;
        frame0.data[1070] = 8'h24; frame0.valid[1070] = 1'b1; frame0.error[1070] = 1'b0;frame0.data[1071] = 8'h25; frame0.valid[1071] = 1'b1; frame0.error[1071] = 1'b0;frame0.data[1072] = 8'h26; frame0.valid[1072] = 1'b1; frame0.error[1072] = 1'b0;frame0.data[1073] = 8'h27; frame0.valid[1073] = 1'b1; frame0.error[1073] = 1'b0;frame0.data[1074] = 8'h28; frame0.valid[1074] = 1'b1; frame0.error[1074] = 1'b0;frame0.data[1075] = 8'h29; frame0.valid[1075] = 1'b1; frame0.error[1075] = 1'b0;frame0.data[1076] = 8'h2A; frame0.valid[1076] = 1'b1; frame0.error[1076] = 1'b0;frame0.data[1077] = 8'h2B; frame0.valid[1077] = 1'b1; frame0.error[1077] = 1'b0;frame0.data[1078] = 8'h2C; frame0.valid[1078] = 1'b1; frame0.error[1078] = 1'b0;frame0.data[1079] = 8'h2D; frame0.valid[1079] = 1'b1; frame0.error[1079] = 1'b0;frame0.data[1080] = 8'h2E; frame0.valid[1080] = 1'b1; frame0.error[1080] = 1'b0;frame0.data[1081] = 8'h2F; frame0.valid[1081] = 1'b1; frame0.error[1081] = 1'b0;frame0.data[1082] = 8'h30; frame0.valid[1082] = 1'b1; frame0.error[1082] = 1'b0;frame0.data[1083] = 8'h31; frame0.valid[1083] = 1'b1; frame0.error[1083] = 1'b0;frame0.data[1084] = 8'h32; frame0.valid[1084] = 1'b1; frame0.error[1084] = 1'b0;frame0.data[1085] = 8'h33; frame0.valid[1085] = 1'b1; frame0.error[1085] = 1'b0;
        frame0.data[1086] = 8'h34; frame0.valid[1086] = 1'b1; frame0.error[1086] = 1'b0;frame0.data[1087] = 8'h35; frame0.valid[1087] = 1'b1; frame0.error[1087] = 1'b0;frame0.data[1088] = 8'h36; frame0.valid[1088] = 1'b1; frame0.error[1088] = 1'b0;frame0.data[1089] = 8'h37; frame0.valid[1089] = 1'b1; frame0.error[1089] = 1'b0;frame0.data[1090] = 8'h38; frame0.valid[1090] = 1'b1; frame0.error[1090] = 1'b0;frame0.data[1091] = 8'h39; frame0.valid[1091] = 1'b1; frame0.error[1091] = 1'b0;frame0.data[1092] = 8'h3A; frame0.valid[1092] = 1'b1; frame0.error[1092] = 1'b0;frame0.data[1093] = 8'h3B; frame0.valid[1093] = 1'b1; frame0.error[1093] = 1'b0;frame0.data[1094] = 8'h3C; frame0.valid[1094] = 1'b1; frame0.error[1094] = 1'b0;frame0.data[1095] = 8'h3D; frame0.valid[1095] = 1'b1; frame0.error[1095] = 1'b0;frame0.data[1096] = 8'h3E; frame0.valid[1096] = 1'b1; frame0.error[1096] = 1'b0;frame0.data[1097] = 8'h3F; frame0.valid[1097] = 1'b1; frame0.error[1097] = 1'b0;frame0.data[1098] = 8'h40; frame0.valid[1098] = 1'b1; frame0.error[1098] = 1'b0;frame0.data[1099] = 8'h41; frame0.valid[1099] = 1'b1; frame0.error[1099] = 1'b0;frame0.data[1100] = 8'h42; frame0.valid[1100] = 1'b1; frame0.error[1100] = 1'b0;frame0.data[1101] = 8'h43; frame0.valid[1101] = 1'b1; frame0.error[1101] = 1'b0;
        frame0.data[1102] = 8'h44; frame0.valid[1102] = 1'b1; frame0.error[1102] = 1'b0;frame0.data[1103] = 8'h45; frame0.valid[1103] = 1'b1; frame0.error[1103] = 1'b0;frame0.data[1104] = 8'h46; frame0.valid[1104] = 1'b1; frame0.error[1104] = 1'b0;frame0.data[1105] = 8'h47; frame0.valid[1105] = 1'b1; frame0.error[1105] = 1'b0;frame0.data[1106] = 8'h48; frame0.valid[1106] = 1'b1; frame0.error[1106] = 1'b0;frame0.data[1107] = 8'h49; frame0.valid[1107] = 1'b1; frame0.error[1107] = 1'b0;frame0.data[1108] = 8'h4A; frame0.valid[1108] = 1'b1; frame0.error[1108] = 1'b0;frame0.data[1109] = 8'h4B; frame0.valid[1109] = 1'b1; frame0.error[1109] = 1'b0;frame0.data[1110] = 8'h4C; frame0.valid[1110] = 1'b1; frame0.error[1110] = 1'b0;frame0.data[1111] = 8'h4D; frame0.valid[1111] = 1'b1; frame0.error[1111] = 1'b0;frame0.data[1112] = 8'h4E; frame0.valid[1112] = 1'b1; frame0.error[1112] = 1'b0;frame0.data[1113] = 8'h4F; frame0.valid[1113] = 1'b1; frame0.error[1113] = 1'b0;frame0.data[1114] = 8'h50; frame0.valid[1114] = 1'b1; frame0.error[1114] = 1'b0;frame0.data[1115] = 8'h51; frame0.valid[1115] = 1'b1; frame0.error[1115] = 1'b0;frame0.data[1116] = 8'h52; frame0.valid[1116] = 1'b1; frame0.error[1116] = 1'b0;frame0.data[1117] = 8'h53; frame0.valid[1117] = 1'b1; frame0.error[1117] = 1'b0;
        frame0.data[1118] = 8'h54; frame0.valid[1118] = 1'b1; frame0.error[1118] = 1'b0;frame0.data[1119] = 8'h55; frame0.valid[1119] = 1'b1; frame0.error[1119] = 1'b0;frame0.data[1120] = 8'h56; frame0.valid[1120] = 1'b1; frame0.error[1120] = 1'b0;frame0.data[1121] = 8'h57; frame0.valid[1121] = 1'b1; frame0.error[1121] = 1'b0;frame0.data[1122] = 8'h58; frame0.valid[1122] = 1'b1; frame0.error[1122] = 1'b0;frame0.data[1123] = 8'h59; frame0.valid[1123] = 1'b1; frame0.error[1123] = 1'b0;frame0.data[1124] = 8'h5A; frame0.valid[1124] = 1'b1; frame0.error[1124] = 1'b0;frame0.data[1125] = 8'h5B; frame0.valid[1125] = 1'b1; frame0.error[1125] = 1'b0;frame0.data[1126] = 8'h5C; frame0.valid[1126] = 1'b1; frame0.error[1126] = 1'b0;frame0.data[1127] = 8'h5D; frame0.valid[1127] = 1'b1; frame0.error[1127] = 1'b0;frame0.data[1128] = 8'h5E; frame0.valid[1128] = 1'b1; frame0.error[1128] = 1'b0;frame0.data[1129] = 8'h5F; frame0.valid[1129] = 1'b1; frame0.error[1129] = 1'b0;frame0.data[1130] = 8'h60; frame0.valid[1130] = 1'b1; frame0.error[1130] = 1'b0;frame0.data[1131] = 8'h61; frame0.valid[1131] = 1'b1; frame0.error[1131] = 1'b0;frame0.data[1132] = 8'h62; frame0.valid[1132] = 1'b1; frame0.error[1132] = 1'b0;frame0.data[1133] = 8'h63; frame0.valid[1133] = 1'b1; frame0.error[1133] = 1'b0;
        frame0.data[1134] = 8'h64; frame0.valid[1134] = 1'b1; frame0.error[1134] = 1'b0;frame0.data[1135] = 8'h65; frame0.valid[1135] = 1'b1; frame0.error[1135] = 1'b0;frame0.data[1136] = 8'h66; frame0.valid[1136] = 1'b1; frame0.error[1136] = 1'b0;frame0.data[1137] = 8'h67; frame0.valid[1137] = 1'b1; frame0.error[1137] = 1'b0;frame0.data[1138] = 8'h68; frame0.valid[1138] = 1'b1; frame0.error[1138] = 1'b0;frame0.data[1139] = 8'h69; frame0.valid[1139] = 1'b1; frame0.error[1139] = 1'b0;frame0.data[1140] = 8'h6A; frame0.valid[1140] = 1'b1; frame0.error[1140] = 1'b0;frame0.data[1141] = 8'h6B; frame0.valid[1141] = 1'b1; frame0.error[1141] = 1'b0;frame0.data[1142] = 8'h6C; frame0.valid[1142] = 1'b1; frame0.error[1142] = 1'b0;frame0.data[1143] = 8'h6D; frame0.valid[1143] = 1'b1; frame0.error[1143] = 1'b0;frame0.data[1144] = 8'h6E; frame0.valid[1144] = 1'b1; frame0.error[1144] = 1'b0;frame0.data[1145] = 8'h6F; frame0.valid[1145] = 1'b1; frame0.error[1145] = 1'b0;frame0.data[1146] = 8'h70; frame0.valid[1146] = 1'b1; frame0.error[1146] = 1'b0;frame0.data[1147] = 8'h71; frame0.valid[1147] = 1'b1; frame0.error[1147] = 1'b0;frame0.data[1148] = 8'h72; frame0.valid[1148] = 1'b1; frame0.error[1148] = 1'b0;frame0.data[1149] = 8'h73; frame0.valid[1149] = 1'b1; frame0.error[1149] = 1'b0;
        frame0.data[1150] = 8'h74; frame0.valid[1150] = 1'b1; frame0.error[1150] = 1'b0;frame0.data[1151] = 8'h75; frame0.valid[1151] = 1'b1; frame0.error[1151] = 1'b0;frame0.data[1152] = 8'h76; frame0.valid[1152] = 1'b1; frame0.error[1152] = 1'b0;frame0.data[1153] = 8'h77; frame0.valid[1153] = 1'b1; frame0.error[1153] = 1'b0;frame0.data[1154] = 8'h78; frame0.valid[1154] = 1'b1; frame0.error[1154] = 1'b0;frame0.data[1155] = 8'h79; frame0.valid[1155] = 1'b1; frame0.error[1155] = 1'b0;frame0.data[1156] = 8'h7A; frame0.valid[1156] = 1'b1; frame0.error[1156] = 1'b0;frame0.data[1157] = 8'h7B; frame0.valid[1157] = 1'b1; frame0.error[1157] = 1'b0;frame0.data[1158] = 8'h7C; frame0.valid[1158] = 1'b1; frame0.error[1158] = 1'b0;frame0.data[1159] = 8'h7D; frame0.valid[1159] = 1'b1; frame0.error[1159] = 1'b0;frame0.data[1160] = 8'h7E; frame0.valid[1160] = 1'b1; frame0.error[1160] = 1'b0;frame0.data[1161] = 8'h7F; frame0.valid[1161] = 1'b1; frame0.error[1161] = 1'b0;frame0.data[1162] = 8'h80; frame0.valid[1162] = 1'b1; frame0.error[1162] = 1'b0;frame0.data[1163] = 8'h81; frame0.valid[1163] = 1'b1; frame0.error[1163] = 1'b0;frame0.data[1164] = 8'h82; frame0.valid[1164] = 1'b1; frame0.error[1164] = 1'b0;frame0.data[1165] = 8'h83; frame0.valid[1165] = 1'b1; frame0.error[1165] = 1'b0;
        frame0.data[1166] = 8'h84; frame0.valid[1166] = 1'b1; frame0.error[1166] = 1'b0;frame0.data[1167] = 8'h85; frame0.valid[1167] = 1'b1; frame0.error[1167] = 1'b0;frame0.data[1168] = 8'h86; frame0.valid[1168] = 1'b1; frame0.error[1168] = 1'b0;frame0.data[1169] = 8'h87; frame0.valid[1169] = 1'b1; frame0.error[1169] = 1'b0;frame0.data[1170] = 8'h88; frame0.valid[1170] = 1'b1; frame0.error[1170] = 1'b0;frame0.data[1171] = 8'h89; frame0.valid[1171] = 1'b1; frame0.error[1171] = 1'b0;frame0.data[1172] = 8'h8A; frame0.valid[1172] = 1'b1; frame0.error[1172] = 1'b0;frame0.data[1173] = 8'h8B; frame0.valid[1173] = 1'b1; frame0.error[1173] = 1'b0;frame0.data[1174] = 8'h8C; frame0.valid[1174] = 1'b1; frame0.error[1174] = 1'b0;frame0.data[1175] = 8'h8D; frame0.valid[1175] = 1'b1; frame0.error[1175] = 1'b0;frame0.data[1176] = 8'h8E; frame0.valid[1176] = 1'b1; frame0.error[1176] = 1'b0;frame0.data[1177] = 8'h8F; frame0.valid[1177] = 1'b1; frame0.error[1177] = 1'b0;frame0.data[1178] = 8'h90; frame0.valid[1178] = 1'b1; frame0.error[1178] = 1'b0;frame0.data[1179] = 8'h91; frame0.valid[1179] = 1'b1; frame0.error[1179] = 1'b0;frame0.data[1180] = 8'h92; frame0.valid[1180] = 1'b1; frame0.error[1180] = 1'b0;frame0.data[1181] = 8'h93; frame0.valid[1181] = 1'b1; frame0.error[1181] = 1'b0;
        frame0.data[1182] = 8'h94; frame0.valid[1182] = 1'b1; frame0.error[1182] = 1'b0;frame0.data[1183] = 8'h95; frame0.valid[1183] = 1'b1; frame0.error[1183] = 1'b0;frame0.data[1184] = 8'h96; frame0.valid[1184] = 1'b1; frame0.error[1184] = 1'b0;frame0.data[1185] = 8'h97; frame0.valid[1185] = 1'b1; frame0.error[1185] = 1'b0;frame0.data[1186] = 8'h98; frame0.valid[1186] = 1'b1; frame0.error[1186] = 1'b0;frame0.data[1187] = 8'h99; frame0.valid[1187] = 1'b1; frame0.error[1187] = 1'b0;frame0.data[1188] = 8'h9A; frame0.valid[1188] = 1'b1; frame0.error[1188] = 1'b0;frame0.data[1189] = 8'h9B; frame0.valid[1189] = 1'b1; frame0.error[1189] = 1'b0;frame0.data[1190] = 8'h9C; frame0.valid[1190] = 1'b1; frame0.error[1190] = 1'b0;frame0.data[1191] = 8'h9D; frame0.valid[1191] = 1'b1; frame0.error[1191] = 1'b0;frame0.data[1192] = 8'h9E; frame0.valid[1192] = 1'b1; frame0.error[1192] = 1'b0;frame0.data[1193] = 8'h9F; frame0.valid[1193] = 1'b1; frame0.error[1193] = 1'b0;frame0.data[1194] = 8'hA0; frame0.valid[1194] = 1'b1; frame0.error[1194] = 1'b0;frame0.data[1195] = 8'hA1; frame0.valid[1195] = 1'b1; frame0.error[1195] = 1'b0;frame0.data[1196] = 8'hA2; frame0.valid[1196] = 1'b1; frame0.error[1196] = 1'b0;frame0.data[1197] = 8'hA3; frame0.valid[1197] = 1'b1; frame0.error[1197] = 1'b0;
        frame0.data[1198] = 8'hA4; frame0.valid[1198] = 1'b1; frame0.error[1198] = 1'b0;frame0.data[1199] = 8'hA5; frame0.valid[1199] = 1'b1; frame0.error[1199] = 1'b0;frame0.data[1200] = 8'hA6; frame0.valid[1200] = 1'b1; frame0.error[1200] = 1'b0;frame0.data[1201] = 8'hA7; frame0.valid[1201] = 1'b1; frame0.error[1201] = 1'b0;frame0.data[1202] = 8'hA8; frame0.valid[1202] = 1'b1; frame0.error[1202] = 1'b0;frame0.data[1203] = 8'hA9; frame0.valid[1203] = 1'b1; frame0.error[1203] = 1'b0;frame0.data[1204] = 8'hAA; frame0.valid[1204] = 1'b1; frame0.error[1204] = 1'b0;frame0.data[1205] = 8'hAB; frame0.valid[1205] = 1'b1; frame0.error[1205] = 1'b0;frame0.data[1206] = 8'hAC; frame0.valid[1206] = 1'b1; frame0.error[1206] = 1'b0;frame0.data[1207] = 8'hAD; frame0.valid[1207] = 1'b1; frame0.error[1207] = 1'b0;frame0.data[1208] = 8'hAE; frame0.valid[1208] = 1'b1; frame0.error[1208] = 1'b0;frame0.data[1209] = 8'hAF; frame0.valid[1209] = 1'b1; frame0.error[1209] = 1'b0;frame0.data[1210] = 8'hB0; frame0.valid[1210] = 1'b1; frame0.error[1210] = 1'b0;frame0.data[1211] = 8'hB1; frame0.valid[1211] = 1'b1; frame0.error[1211] = 1'b0;frame0.data[1212] = 8'hB2; frame0.valid[1212] = 1'b1; frame0.error[1212] = 1'b0;frame0.data[1213] = 8'hB3; frame0.valid[1213] = 1'b1; frame0.error[1213] = 1'b0;
        frame0.data[1214] = 8'hB4; frame0.valid[1214] = 1'b1; frame0.error[1214] = 1'b0;frame0.data[1215] = 8'hB5; frame0.valid[1215] = 1'b1; frame0.error[1215] = 1'b0;frame0.data[1216] = 8'hB6; frame0.valid[1216] = 1'b1; frame0.error[1216] = 1'b0;frame0.data[1217] = 8'hB7; frame0.valid[1217] = 1'b1; frame0.error[1217] = 1'b0;frame0.data[1218] = 8'hB8; frame0.valid[1218] = 1'b1; frame0.error[1218] = 1'b0;frame0.data[1219] = 8'hB9; frame0.valid[1219] = 1'b1; frame0.error[1219] = 1'b0;frame0.data[1220] = 8'hBA; frame0.valid[1220] = 1'b1; frame0.error[1220] = 1'b0;frame0.data[1221] = 8'hBB; frame0.valid[1221] = 1'b1; frame0.error[1221] = 1'b0;frame0.data[1222] = 8'hBC; frame0.valid[1222] = 1'b1; frame0.error[1222] = 1'b0;frame0.data[1223] = 8'hBD; frame0.valid[1223] = 1'b1; frame0.error[1223] = 1'b0;frame0.data[1224] = 8'hBE; frame0.valid[1224] = 1'b1; frame0.error[1224] = 1'b0;frame0.data[1225] = 8'hBF; frame0.valid[1225] = 1'b1; frame0.error[1225] = 1'b0;frame0.data[1226] = 8'hC0; frame0.valid[1226] = 1'b1; frame0.error[1226] = 1'b0;frame0.data[1227] = 8'hC1; frame0.valid[1227] = 1'b1; frame0.error[1227] = 1'b0;frame0.data[1228] = 8'hC2; frame0.valid[1228] = 1'b1; frame0.error[1228] = 1'b0;frame0.data[1229] = 8'hC3; frame0.valid[1229] = 1'b1; frame0.error[1229] = 1'b0;
        frame0.data[1230] = 8'hC4; frame0.valid[1230] = 1'b1; frame0.error[1230] = 1'b0;frame0.data[1231] = 8'hC5; frame0.valid[1231] = 1'b1; frame0.error[1231] = 1'b0;frame0.data[1232] = 8'hC6; frame0.valid[1232] = 1'b1; frame0.error[1232] = 1'b0;frame0.data[1233] = 8'hC7; frame0.valid[1233] = 1'b1; frame0.error[1233] = 1'b0;frame0.data[1234] = 8'hC8; frame0.valid[1234] = 1'b1; frame0.error[1234] = 1'b0;frame0.data[1235] = 8'hC9; frame0.valid[1235] = 1'b1; frame0.error[1235] = 1'b0;frame0.data[1236] = 8'hCA; frame0.valid[1236] = 1'b1; frame0.error[1236] = 1'b0;frame0.data[1237] = 8'hCB; frame0.valid[1237] = 1'b1; frame0.error[1237] = 1'b0;frame0.data[1238] = 8'hCC; frame0.valid[1238] = 1'b1; frame0.error[1238] = 1'b0;frame0.data[1239] = 8'hCD; frame0.valid[1239] = 1'b1; frame0.error[1239] = 1'b0;frame0.data[1240] = 8'hCE; frame0.valid[1240] = 1'b1; frame0.error[1240] = 1'b0;frame0.data[1241] = 8'hCF; frame0.valid[1241] = 1'b1; frame0.error[1241] = 1'b0;frame0.data[1242] = 8'hD0; frame0.valid[1242] = 1'b1; frame0.error[1242] = 1'b0;frame0.data[1243] = 8'hD1; frame0.valid[1243] = 1'b1; frame0.error[1243] = 1'b0;frame0.data[1244] = 8'hD2; frame0.valid[1244] = 1'b1; frame0.error[1244] = 1'b0;frame0.data[1245] = 8'hD3; frame0.valid[1245] = 1'b1; frame0.error[1245] = 1'b0;
        frame0.data[1246] = 8'hD4; frame0.valid[1246] = 1'b1; frame0.error[1246] = 1'b0;frame0.data[1247] = 8'hD5; frame0.valid[1247] = 1'b1; frame0.error[1247] = 1'b0;frame0.data[1248] = 8'hD6; frame0.valid[1248] = 1'b1; frame0.error[1248] = 1'b0;frame0.data[1249] = 8'hD7; frame0.valid[1249] = 1'b1; frame0.error[1249] = 1'b0;frame0.data[1250] = 8'hD8; frame0.valid[1250] = 1'b1; frame0.error[1250] = 1'b0;frame0.data[1251] = 8'hD9; frame0.valid[1251] = 1'b1; frame0.error[1251] = 1'b0;frame0.data[1252] = 8'hDA; frame0.valid[1252] = 1'b1; frame0.error[1252] = 1'b0;frame0.data[1253] = 8'hDB; frame0.valid[1253] = 1'b1; frame0.error[1253] = 1'b0;frame0.data[1254] = 8'hDC; frame0.valid[1254] = 1'b1; frame0.error[1254] = 1'b0;frame0.data[1255] = 8'hDD; frame0.valid[1255] = 1'b1; frame0.error[1255] = 1'b0;frame0.data[1256] = 8'hDE; frame0.valid[1256] = 1'b1; frame0.error[1256] = 1'b0;frame0.data[1257] = 8'hDF; frame0.valid[1257] = 1'b1; frame0.error[1257] = 1'b0;frame0.data[1258] = 8'hE0; frame0.valid[1258] = 1'b1; frame0.error[1258] = 1'b0;frame0.data[1259] = 8'hE1; frame0.valid[1259] = 1'b1; frame0.error[1259] = 1'b0;frame0.data[1260] = 8'hE2; frame0.valid[1260] = 1'b1; frame0.error[1260] = 1'b0;frame0.data[1261] = 8'hE3; frame0.valid[1261] = 1'b1; frame0.error[1261] = 1'b0;
        frame0.data[1262] = 8'hE4; frame0.valid[1262] = 1'b1; frame0.error[1262] = 1'b0;frame0.data[1263] = 8'hE5; frame0.valid[1263] = 1'b1; frame0.error[1263] = 1'b0;frame0.data[1264] = 8'hE6; frame0.valid[1264] = 1'b1; frame0.error[1264] = 1'b0;frame0.data[1265] = 8'hE7; frame0.valid[1265] = 1'b1; frame0.error[1265] = 1'b0;frame0.data[1266] = 8'hE8; frame0.valid[1266] = 1'b1; frame0.error[1266] = 1'b0;frame0.data[1267] = 8'hE9; frame0.valid[1267] = 1'b1; frame0.error[1267] = 1'b0;frame0.data[1268] = 8'hEA; frame0.valid[1268] = 1'b1; frame0.error[1268] = 1'b0;frame0.data[1269] = 8'hEB; frame0.valid[1269] = 1'b1; frame0.error[1269] = 1'b0;frame0.data[1270] = 8'hEC; frame0.valid[1270] = 1'b1; frame0.error[1270] = 1'b0;frame0.data[1271] = 8'hED; frame0.valid[1271] = 1'b1; frame0.error[1271] = 1'b0;frame0.data[1272] = 8'hEE; frame0.valid[1272] = 1'b1; frame0.error[1272] = 1'b0;frame0.data[1273] = 8'hEF; frame0.valid[1273] = 1'b1; frame0.error[1273] = 1'b0;frame0.data[1274] = 8'hF0; frame0.valid[1274] = 1'b1; frame0.error[1274] = 1'b0;frame0.data[1275] = 8'hF1; frame0.valid[1275] = 1'b1; frame0.error[1275] = 1'b0;frame0.data[1276] = 8'hF2; frame0.valid[1276] = 1'b1; frame0.error[1276] = 1'b0;frame0.data[1277] = 8'hF3; frame0.valid[1277] = 1'b1; frame0.error[1277] = 1'b0;
        frame0.data[1278] = 8'hF4; frame0.valid[1278] = 1'b1; frame0.error[1278] = 1'b0;frame0.data[1279] = 8'hF5; frame0.valid[1279] = 1'b1; frame0.error[1279] = 1'b0;frame0.data[1280] = 8'hF6; frame0.valid[1280] = 1'b1; frame0.error[1280] = 1'b0;frame0.data[1281] = 8'hF7; frame0.valid[1281] = 1'b1; frame0.error[1281] = 1'b0;frame0.data[1282] = 8'hF8; frame0.valid[1282] = 1'b1; frame0.error[1282] = 1'b0;frame0.data[1283] = 8'hF9; frame0.valid[1283] = 1'b1; frame0.error[1283] = 1'b0;frame0.data[1284] = 8'hFA; frame0.valid[1284] = 1'b1; frame0.error[1284] = 1'b0;frame0.data[1285] = 8'hFB; frame0.valid[1285] = 1'b1; frame0.error[1285] = 1'b0;frame0.data[1286] = 8'hFC; frame0.valid[1286] = 1'b1; frame0.error[1286] = 1'b0;frame0.data[1287] = 8'hFD; frame0.valid[1287] = 1'b1; frame0.error[1287] = 1'b0;frame0.data[1288] = 8'hFE; frame0.valid[1288] = 1'b1; frame0.error[1288] = 1'b0;frame0.data[1289] = 8'h00; frame0.valid[1289] = 1'b1; frame0.error[1289] = 1'b0;frame0.data[1290] = 8'h01; frame0.valid[1290] = 1'b1; frame0.error[1290] = 1'b0;frame0.data[1291] = 8'h02; frame0.valid[1291] = 1'b1; frame0.error[1291] = 1'b0;frame0.data[1292] = 8'h03; frame0.valid[1292] = 1'b1; frame0.error[1292] = 1'b0;frame0.data[1293] = 8'h04; frame0.valid[1293] = 1'b1; frame0.error[1293] = 1'b0;
        frame0.data[1294] = 8'h05; frame0.valid[1294] = 1'b1; frame0.error[1294] = 1'b0;frame0.data[1295] = 8'h06; frame0.valid[1295] = 1'b1; frame0.error[1295] = 1'b0;frame0.data[1296] = 8'h07; frame0.valid[1296] = 1'b1; frame0.error[1296] = 1'b0;frame0.data[1297] = 8'h08; frame0.valid[1297] = 1'b1; frame0.error[1297] = 1'b0;frame0.data[1298] = 8'h09; frame0.valid[1298] = 1'b1; frame0.error[1298] = 1'b0;frame0.data[1299] = 8'h0A; frame0.valid[1299] = 1'b1; frame0.error[1299] = 1'b0;frame0.data[1300] = 8'h0B; frame0.valid[1300] = 1'b1; frame0.error[1300] = 1'b0;frame0.data[1301] = 8'h0C; frame0.valid[1301] = 1'b1; frame0.error[1301] = 1'b0;frame0.data[1302] = 8'h0D; frame0.valid[1302] = 1'b1; frame0.error[1302] = 1'b0;frame0.data[1303] = 8'h0E; frame0.valid[1303] = 1'b1; frame0.error[1303] = 1'b0;frame0.data[1304] = 8'h0F; frame0.valid[1304] = 1'b1; frame0.error[1304] = 1'b0;frame0.data[1305] = 8'h10; frame0.valid[1305] = 1'b1; frame0.error[1305] = 1'b0;frame0.data[1306] = 8'h11; frame0.valid[1306] = 1'b1; frame0.error[1306] = 1'b0;frame0.data[1307] = 8'h12; frame0.valid[1307] = 1'b1; frame0.error[1307] = 1'b0;frame0.data[1308] = 8'h13; frame0.valid[1308] = 1'b1; frame0.error[1308] = 1'b0;frame0.data[1309] = 8'h14; frame0.valid[1309] = 1'b1; frame0.error[1309] = 1'b0;
        frame0.data[1310] = 8'h15; frame0.valid[1310] = 1'b1; frame0.error[1310] = 1'b0;frame0.data[1311] = 8'h16; frame0.valid[1311] = 1'b1; frame0.error[1311] = 1'b0;frame0.data[1312] = 8'h17; frame0.valid[1312] = 1'b1; frame0.error[1312] = 1'b0;frame0.data[1313] = 8'h18; frame0.valid[1313] = 1'b1; frame0.error[1313] = 1'b0;frame0.data[1314] = 8'h19; frame0.valid[1314] = 1'b1; frame0.error[1314] = 1'b0;frame0.data[1315] = 8'h1A; frame0.valid[1315] = 1'b1; frame0.error[1315] = 1'b0;frame0.data[1316] = 8'h1B; frame0.valid[1316] = 1'b1; frame0.error[1316] = 1'b0;frame0.data[1317] = 8'h1C; frame0.valid[1317] = 1'b1; frame0.error[1317] = 1'b0;frame0.data[1318] = 8'h1D; frame0.valid[1318] = 1'b1; frame0.error[1318] = 1'b0;frame0.data[1319] = 8'h1E; frame0.valid[1319] = 1'b1; frame0.error[1319] = 1'b0;frame0.data[1320] = 8'h1F; frame0.valid[1320] = 1'b1; frame0.error[1320] = 1'b0;frame0.data[1321] = 8'h20; frame0.valid[1321] = 1'b1; frame0.error[1321] = 1'b0;frame0.data[1322] = 8'h21; frame0.valid[1322] = 1'b1; frame0.error[1322] = 1'b0;frame0.data[1323] = 8'h22; frame0.valid[1323] = 1'b1; frame0.error[1323] = 1'b0;frame0.data[1324] = 8'h23; frame0.valid[1324] = 1'b1; frame0.error[1324] = 1'b0;frame0.data[1325] = 8'h24; frame0.valid[1325] = 1'b1; frame0.error[1325] = 1'b0;
        frame0.data[1326] = 8'h25; frame0.valid[1326] = 1'b1; frame0.error[1326] = 1'b0;frame0.data[1327] = 8'h26; frame0.valid[1327] = 1'b1; frame0.error[1327] = 1'b0;frame0.data[1328] = 8'h27; frame0.valid[1328] = 1'b1; frame0.error[1328] = 1'b0;frame0.data[1329] = 8'h28; frame0.valid[1329] = 1'b1; frame0.error[1329] = 1'b0;frame0.data[1330] = 8'h29; frame0.valid[1330] = 1'b1; frame0.error[1330] = 1'b0;frame0.data[1331] = 8'h2A; frame0.valid[1331] = 1'b1; frame0.error[1331] = 1'b0;frame0.data[1332] = 8'h2B; frame0.valid[1332] = 1'b1; frame0.error[1332] = 1'b0;frame0.data[1333] = 8'h2C; frame0.valid[1333] = 1'b1; frame0.error[1333] = 1'b0;frame0.data[1334] = 8'h2D; frame0.valid[1334] = 1'b1; frame0.error[1334] = 1'b0;frame0.data[1335] = 8'h2E; frame0.valid[1335] = 1'b1; frame0.error[1335] = 1'b0;frame0.data[1336] = 8'h2F; frame0.valid[1336] = 1'b1; frame0.error[1336] = 1'b0;frame0.data[1337] = 8'h30; frame0.valid[1337] = 1'b1; frame0.error[1337] = 1'b0;frame0.data[1338] = 8'h31; frame0.valid[1338] = 1'b1; frame0.error[1338] = 1'b0;frame0.data[1339] = 8'h32; frame0.valid[1339] = 1'b1; frame0.error[1339] = 1'b0;frame0.data[1340] = 8'h33; frame0.valid[1340] = 1'b1; frame0.error[1340] = 1'b0;frame0.data[1341] = 8'h34; frame0.valid[1341] = 1'b1; frame0.error[1341] = 1'b0;
        frame0.data[1342] = 8'h35; frame0.valid[1342] = 1'b1; frame0.error[1342] = 1'b0;frame0.data[1343] = 8'h36; frame0.valid[1343] = 1'b1; frame0.error[1343] = 1'b0;frame0.data[1344] = 8'h37; frame0.valid[1344] = 1'b1; frame0.error[1344] = 1'b0;frame0.data[1345] = 8'h38; frame0.valid[1345] = 1'b1; frame0.error[1345] = 1'b0;frame0.data[1346] = 8'h39; frame0.valid[1346] = 1'b1; frame0.error[1346] = 1'b0;frame0.data[1347] = 8'h3A; frame0.valid[1347] = 1'b1; frame0.error[1347] = 1'b0;frame0.data[1348] = 8'h3B; frame0.valid[1348] = 1'b1; frame0.error[1348] = 1'b0;frame0.data[1349] = 8'h3C; frame0.valid[1349] = 1'b1; frame0.error[1349] = 1'b0;frame0.data[1350] = 8'h3D; frame0.valid[1350] = 1'b1; frame0.error[1350] = 1'b0;frame0.data[1351] = 8'h3E; frame0.valid[1351] = 1'b1; frame0.error[1351] = 1'b0;frame0.data[1352] = 8'h3F; frame0.valid[1352] = 1'b1; frame0.error[1352] = 1'b0;frame0.data[1353] = 8'h40; frame0.valid[1353] = 1'b1; frame0.error[1353] = 1'b0;frame0.data[1354] = 8'h41; frame0.valid[1354] = 1'b1; frame0.error[1354] = 1'b0;frame0.data[1355] = 8'h42; frame0.valid[1355] = 1'b1; frame0.error[1355] = 1'b0;frame0.data[1356] = 8'h43; frame0.valid[1356] = 1'b1; frame0.error[1356] = 1'b0;frame0.data[1357] = 8'h44; frame0.valid[1357] = 1'b1; frame0.error[1357] = 1'b0;
        frame0.data[1358] = 8'h45; frame0.valid[1358] = 1'b1; frame0.error[1358] = 1'b0;frame0.data[1359] = 8'h46; frame0.valid[1359] = 1'b1; frame0.error[1359] = 1'b0;frame0.data[1360] = 8'h47; frame0.valid[1360] = 1'b1; frame0.error[1360] = 1'b0;frame0.data[1361] = 8'h48; frame0.valid[1361] = 1'b1; frame0.error[1361] = 1'b0;frame0.data[1362] = 8'h49; frame0.valid[1362] = 1'b1; frame0.error[1362] = 1'b0;frame0.data[1363] = 8'h4A; frame0.valid[1363] = 1'b1; frame0.error[1363] = 1'b0;frame0.data[1364] = 8'h4B; frame0.valid[1364] = 1'b1; frame0.error[1364] = 1'b0;frame0.data[1365] = 8'h4C; frame0.valid[1365] = 1'b1; frame0.error[1365] = 1'b0;frame0.data[1366] = 8'h4D; frame0.valid[1366] = 1'b1; frame0.error[1366] = 1'b0;frame0.data[1367] = 8'h4E; frame0.valid[1367] = 1'b1; frame0.error[1367] = 1'b0;frame0.data[1368] = 8'h4F; frame0.valid[1368] = 1'b1; frame0.error[1368] = 1'b0;frame0.data[1369] = 8'h50; frame0.valid[1369] = 1'b1; frame0.error[1369] = 1'b0;frame0.data[1370] = 8'h51; frame0.valid[1370] = 1'b1; frame0.error[1370] = 1'b0;frame0.data[1371] = 8'h52; frame0.valid[1371] = 1'b1; frame0.error[1371] = 1'b0;frame0.data[1372] = 8'h53; frame0.valid[1372] = 1'b1; frame0.error[1372] = 1'b0;frame0.data[1373] = 8'h54; frame0.valid[1373] = 1'b1; frame0.error[1373] = 1'b0;
        frame0.data[1374] = 8'h55; frame0.valid[1374] = 1'b1; frame0.error[1374] = 1'b0;frame0.data[1375] = 8'h56; frame0.valid[1375] = 1'b1; frame0.error[1375] = 1'b0;frame0.data[1376] = 8'h57; frame0.valid[1376] = 1'b1; frame0.error[1376] = 1'b0;frame0.data[1377] = 8'h58; frame0.valid[1377] = 1'b1; frame0.error[1377] = 1'b0;frame0.data[1378] = 8'h59; frame0.valid[1378] = 1'b1; frame0.error[1378] = 1'b0;frame0.data[1379] = 8'h5A; frame0.valid[1379] = 1'b1; frame0.error[1379] = 1'b0;frame0.data[1380] = 8'h5B; frame0.valid[1380] = 1'b1; frame0.error[1380] = 1'b0;frame0.data[1381] = 8'h5C; frame0.valid[1381] = 1'b1; frame0.error[1381] = 1'b0;frame0.data[1382] = 8'h5D; frame0.valid[1382] = 1'b1; frame0.error[1382] = 1'b0;frame0.data[1383] = 8'h5E; frame0.valid[1383] = 1'b1; frame0.error[1383] = 1'b0;frame0.data[1384] = 8'h5F; frame0.valid[1384] = 1'b1; frame0.error[1384] = 1'b0;frame0.data[1385] = 8'h60; frame0.valid[1385] = 1'b1; frame0.error[1385] = 1'b0;frame0.data[1386] = 8'h61; frame0.valid[1386] = 1'b1; frame0.error[1386] = 1'b0;frame0.data[1387] = 8'h62; frame0.valid[1387] = 1'b1; frame0.error[1387] = 1'b0;frame0.data[1388] = 8'h63; frame0.valid[1388] = 1'b1; frame0.error[1388] = 1'b0;frame0.data[1389] = 8'h64; frame0.valid[1389] = 1'b1; frame0.error[1389] = 1'b0;
        frame0.data[1390] = 8'h65; frame0.valid[1390] = 1'b1; frame0.error[1390] = 1'b0;frame0.data[1391] = 8'h66; frame0.valid[1391] = 1'b1; frame0.error[1391] = 1'b0;frame0.data[1392] = 8'h67; frame0.valid[1392] = 1'b1; frame0.error[1392] = 1'b0;frame0.data[1393] = 8'h68; frame0.valid[1393] = 1'b1; frame0.error[1393] = 1'b0;frame0.data[1394] = 8'h69; frame0.valid[1394] = 1'b1; frame0.error[1394] = 1'b0;frame0.data[1395] = 8'h6A; frame0.valid[1395] = 1'b1; frame0.error[1395] = 1'b0;frame0.data[1396] = 8'h6B; frame0.valid[1396] = 1'b1; frame0.error[1396] = 1'b0;frame0.data[1397] = 8'h6C; frame0.valid[1397] = 1'b1; frame0.error[1397] = 1'b0;frame0.data[1398] = 8'h6D; frame0.valid[1398] = 1'b1; frame0.error[1398] = 1'b0;frame0.data[1399] = 8'h6E; frame0.valid[1399] = 1'b1; frame0.error[1399] = 1'b0;frame0.data[1400] = 8'h6F; frame0.valid[1400] = 1'b1; frame0.error[1400] = 1'b0;frame0.data[1401] = 8'h70; frame0.valid[1401] = 1'b1; frame0.error[1401] = 1'b0;frame0.data[1402] = 8'h71; frame0.valid[1402] = 1'b1; frame0.error[1402] = 1'b0;frame0.data[1403] = 8'h72; frame0.valid[1403] = 1'b1; frame0.error[1403] = 1'b0;frame0.data[1404] = 8'h73; frame0.valid[1404] = 1'b1; frame0.error[1404] = 1'b0;frame0.data[1405] = 8'h74; frame0.valid[1405] = 1'b1; frame0.error[1405] = 1'b0;
        frame0.data[1406] = 8'h75; frame0.valid[1406] = 1'b1; frame0.error[1406] = 1'b0;frame0.data[1407] = 8'h76; frame0.valid[1407] = 1'b1; frame0.error[1407] = 1'b0;frame0.data[1408] = 8'h77; frame0.valid[1408] = 1'b1; frame0.error[1408] = 1'b0;frame0.data[1409] = 8'h78; frame0.valid[1409] = 1'b1; frame0.error[1409] = 1'b0;frame0.data[1410] = 8'h79; frame0.valid[1410] = 1'b1; frame0.error[1410] = 1'b0;frame0.data[1411] = 8'h7A; frame0.valid[1411] = 1'b1; frame0.error[1411] = 1'b0;frame0.data[1412] = 8'h7B; frame0.valid[1412] = 1'b1; frame0.error[1412] = 1'b0;frame0.data[1413] = 8'h7C; frame0.valid[1413] = 1'b1; frame0.error[1413] = 1'b0;frame0.data[1414] = 8'h7D; frame0.valid[1414] = 1'b1; frame0.error[1414] = 1'b0;frame0.data[1415] = 8'h7E; frame0.valid[1415] = 1'b1; frame0.error[1415] = 1'b0;frame0.data[1416] = 8'h7F; frame0.valid[1416] = 1'b1; frame0.error[1416] = 1'b0;frame0.data[1417] = 8'h80; frame0.valid[1417] = 1'b1; frame0.error[1417] = 1'b0;frame0.data[1418] = 8'h81; frame0.valid[1418] = 1'b1; frame0.error[1418] = 1'b0;frame0.data[1419] = 8'h82; frame0.valid[1419] = 1'b1; frame0.error[1419] = 1'b0;frame0.data[1420] = 8'h83; frame0.valid[1420] = 1'b1; frame0.error[1420] = 1'b0;frame0.data[1421] = 8'h84; frame0.valid[1421] = 1'b1; frame0.error[1421] = 1'b0;
        frame0.data[1422] = 8'h85; frame0.valid[1422] = 1'b1; frame0.error[1422] = 1'b0;frame0.data[1423] = 8'h86; frame0.valid[1423] = 1'b1; frame0.error[1423] = 1'b0;frame0.data[1424] = 8'h87; frame0.valid[1424] = 1'b1; frame0.error[1424] = 1'b0;frame0.data[1425] = 8'h88; frame0.valid[1425] = 1'b1; frame0.error[1425] = 1'b0;frame0.data[1426] = 8'h89; frame0.valid[1426] = 1'b1; frame0.error[1426] = 1'b0;frame0.data[1427] = 8'h8A; frame0.valid[1427] = 1'b1; frame0.error[1427] = 1'b0;frame0.data[1428] = 8'h8B; frame0.valid[1428] = 1'b1; frame0.error[1428] = 1'b0;frame0.data[1429] = 8'h8C; frame0.valid[1429] = 1'b1; frame0.error[1429] = 1'b0;frame0.data[1430] = 8'h8D; frame0.valid[1430] = 1'b1; frame0.error[1430] = 1'b0;frame0.data[1431] = 8'h8E; frame0.valid[1431] = 1'b1; frame0.error[1431] = 1'b0;frame0.data[1432] = 8'h8F; frame0.valid[1432] = 1'b1; frame0.error[1432] = 1'b0;frame0.data[1433] = 8'h90; frame0.valid[1433] = 1'b1; frame0.error[1433] = 1'b0;frame0.data[1434] = 8'h91; frame0.valid[1434] = 1'b1; frame0.error[1434] = 1'b0;frame0.data[1435] = 8'h92; frame0.valid[1435] = 1'b1; frame0.error[1435] = 1'b0;frame0.data[1436] = 8'h93; frame0.valid[1436] = 1'b1; frame0.error[1436] = 1'b0;frame0.data[1437] = 8'h94; frame0.valid[1437] = 1'b1; frame0.error[1437] = 1'b0;
        frame0.data[1438] = 8'h95; frame0.valid[1438] = 1'b1; frame0.error[1438] = 1'b0;frame0.data[1439] = 8'h96; frame0.valid[1439] = 1'b1; frame0.error[1439] = 1'b0;frame0.data[1440] = 8'h97; frame0.valid[1440] = 1'b1; frame0.error[1440] = 1'b0;frame0.data[1441] = 8'h98; frame0.valid[1441] = 1'b1; frame0.error[1441] = 1'b0;frame0.data[1442] = 8'h99; frame0.valid[1442] = 1'b1; frame0.error[1442] = 1'b0;frame0.data[1443] = 8'h9A; frame0.valid[1443] = 1'b1; frame0.error[1443] = 1'b0;frame0.data[1444] = 8'h9B; frame0.valid[1444] = 1'b1; frame0.error[1444] = 1'b0;frame0.data[1445] = 8'h9C; frame0.valid[1445] = 1'b1; frame0.error[1445] = 1'b0;frame0.data[1446] = 8'h9D; frame0.valid[1446] = 1'b1; frame0.error[1446] = 1'b0;frame0.data[1447] = 8'h9E; frame0.valid[1447] = 1'b1; frame0.error[1447] = 1'b0;frame0.data[1448] = 8'h9F; frame0.valid[1448] = 1'b1; frame0.error[1448] = 1'b0;frame0.data[1449] = 8'hA0; frame0.valid[1449] = 1'b1; frame0.error[1449] = 1'b0;frame0.data[1450] = 8'hA1; frame0.valid[1450] = 1'b1; frame0.error[1450] = 1'b0;frame0.data[1451] = 8'hA2; frame0.valid[1451] = 1'b1; frame0.error[1451] = 1'b0;frame0.data[1452] = 8'hA3; frame0.valid[1452] = 1'b1; frame0.error[1452] = 1'b0;frame0.data[1453] = 8'hA4; frame0.valid[1453] = 1'b1; frame0.error[1453] = 1'b0;
        frame0.data[1454] = 8'hA5; frame0.valid[1454] = 1'b1; frame0.error[1454] = 1'b0;frame0.data[1455] = 8'hA6; frame0.valid[1455] = 1'b1; frame0.error[1455] = 1'b0;frame0.data[1456] = 8'hA7; frame0.valid[1456] = 1'b1; frame0.error[1456] = 1'b0;frame0.data[1457] = 8'hA8; frame0.valid[1457] = 1'b1; frame0.error[1457] = 1'b0;frame0.data[1458] = 8'hA9; frame0.valid[1458] = 1'b1; frame0.error[1458] = 1'b0;frame0.data[1459] = 8'hAA; frame0.valid[1459] = 1'b1; frame0.error[1459] = 1'b0;frame0.data[1460] = 8'hAB; frame0.valid[1460] = 1'b1; frame0.error[1460] = 1'b0;frame0.data[1461] = 8'hAC; frame0.valid[1461] = 1'b1; frame0.error[1461] = 1'b0;frame0.data[1462] = 8'hAD; frame0.valid[1462] = 1'b1; frame0.error[1462] = 1'b0;frame0.data[1463] = 8'hAE; frame0.valid[1463] = 1'b1; frame0.error[1463] = 1'b0;frame0.data[1464] = 8'hAF; frame0.valid[1464] = 1'b1; frame0.error[1464] = 1'b0;frame0.data[1465] = 8'hB0; frame0.valid[1465] = 1'b1; frame0.error[1465] = 1'b0;frame0.data[1466] = 8'hB1; frame0.valid[1466] = 1'b1; frame0.error[1466] = 1'b0;frame0.data[1467] = 8'hB2; frame0.valid[1467] = 1'b1; frame0.error[1467] = 1'b0;frame0.data[1468] = 8'hB3; frame0.valid[1468] = 1'b1; frame0.error[1468] = 1'b0;frame0.data[1469] = 8'hB4; frame0.valid[1469] = 1'b1; frame0.error[1469] = 1'b0;
        frame0.data[1470] = 8'hB5; frame0.valid[1470] = 1'b1; frame0.error[1470] = 1'b0;frame0.data[1471] = 8'hB6; frame0.valid[1471] = 1'b1; frame0.error[1471] = 1'b0;frame0.data[1472] = 8'hB7; frame0.valid[1472] = 1'b1; frame0.error[1472] = 1'b0;frame0.data[1473] = 8'hB8; frame0.valid[1473] = 1'b1; frame0.error[1473] = 1'b0;frame0.data[1474] = 8'hB9; frame0.valid[1474] = 1'b1; frame0.error[1474] = 1'b0;frame0.data[1475] = 8'hBA; frame0.valid[1475] = 1'b1; frame0.error[1475] = 1'b0;frame0.data[1476] = 8'hBB; frame0.valid[1476] = 1'b1; frame0.error[1476] = 1'b0;frame0.data[1477] = 8'hBC; frame0.valid[1477] = 1'b1; frame0.error[1477] = 1'b0;frame0.data[1478] = 8'hBD; frame0.valid[1478] = 1'b1; frame0.error[1478] = 1'b0;frame0.data[1479] = 8'hBE; frame0.valid[1479] = 1'b1; frame0.error[1479] = 1'b0;frame0.data[1480] = 8'hBF; frame0.valid[1480] = 1'b1; frame0.error[1480] = 1'b0;frame0.data[1481] = 8'hC0; frame0.valid[1481] = 1'b1; frame0.error[1481] = 1'b0;frame0.data[1482] = 8'hC1; frame0.valid[1482] = 1'b1; frame0.error[1482] = 1'b0;frame0.data[1483] = 8'hC2; frame0.valid[1483] = 1'b1; frame0.error[1483] = 1'b0;frame0.data[1484] = 8'hC3; frame0.valid[1484] = 1'b1; frame0.error[1484] = 1'b0;frame0.data[1485] = 8'hC4; frame0.valid[1485] = 1'b1; frame0.error[1485] = 1'b0;
        frame0.data[1486] = 8'hC5; frame0.valid[1486] = 1'b1; frame0.error[1486] = 1'b0;frame0.data[1487] = 8'hC6; frame0.valid[1487] = 1'b1; frame0.error[1487] = 1'b0;frame0.data[1488] = 8'hC7; frame0.valid[1488] = 1'b1; frame0.error[1488] = 1'b0;frame0.data[1489] = 8'hC8; frame0.valid[1489] = 1'b1; frame0.error[1489] = 1'b0;frame0.data[1490] = 8'hC9; frame0.valid[1490] = 1'b1; frame0.error[1490] = 1'b0;frame0.data[1491] = 8'hCA; frame0.valid[1491] = 1'b1; frame0.error[1491] = 1'b0;frame0.data[1492] = 8'hCB; frame0.valid[1492] = 1'b1; frame0.error[1492] = 1'b0;frame0.data[1493] = 8'hCC; frame0.valid[1493] = 1'b1; frame0.error[1493] = 1'b0;frame0.data[1494] = 8'hCD; frame0.valid[1494] = 1'b1; frame0.error[1494] = 1'b0;frame0.data[1495] = 8'hCE; frame0.valid[1495] = 1'b1; frame0.error[1495] = 1'b0;frame0.data[1496] = 8'hCF; frame0.valid[1496] = 1'b1; frame0.error[1496] = 1'b0;frame0.data[1497] = 8'hD0; frame0.valid[1497] = 1'b1; frame0.error[1497] = 1'b0;frame0.data[1498] = 8'hD1; frame0.valid[1498] = 1'b1; frame0.error[1498] = 1'b0;frame0.data[1499] = 8'hD2; frame0.valid[1499] = 1'b1; frame0.error[1499] = 1'b0;frame0.data[1500] = 8'hD3; frame0.valid[1500] = 1'b1; frame0.error[1500] = 1'b0;frame0.data[1501] = 8'hD4; frame0.valid[1501] = 1'b1; frame0.error[1501] = 1'b0;
        frame0.data[1502] = 8'hD5; frame0.valid[1502] = 1'b1; frame0.error[1502] = 1'b0;frame0.data[1503] = 8'hD6; frame0.valid[1503] = 1'b1; frame0.error[1503] = 1'b0;frame0.data[1504] = 8'hD7; frame0.valid[1504] = 1'b1; frame0.error[1504] = 1'b0;frame0.data[1505] = 8'hD8; frame0.valid[1505] = 1'b1; frame0.error[1505] = 1'b0;frame0.data[1506] = 8'hD9; frame0.valid[1506] = 1'b1; frame0.error[1506] = 1'b0;frame0.data[1507] = 8'hDA; frame0.valid[1507] = 1'b1; frame0.error[1507] = 1'b0;frame0.data[1508] = 8'hDB; frame0.valid[1508] = 1'b1; frame0.error[1508] = 1'b0;frame0.data[1509] = 8'hDC; frame0.valid[1509] = 1'b1; frame0.error[1509] = 1'b0;frame0.data[1510] = 8'hDD; frame0.valid[1510] = 1'b1; frame0.error[1510] = 1'b0;frame0.data[1511] = 8'hDE; frame0.valid[1511] = 1'b1; frame0.error[1511] = 1'b0;frame0.data[1512] = 8'hDF; frame0.valid[1512] = 1'b1; frame0.error[1512] = 1'b0;frame0.data[1513] = 8'hE0; frame0.valid[1513] = 1'b1; frame0.error[1513] = 1'b0;
        // unused
        frame0.data[1514] = 8'h00;  frame0.valid[1514] = 1'b0;  frame0.error[1514] = 1'b0;
        frame0.data[1515] = 8'h00;  frame0.valid[1515] = 1'b0;  frame0.error[1515] = 1'b0;

        // No error in this frame
        frame0.bad_frame  = 1'b0;

        //-----------
        // Frame 1
        // PTP message
        //-----------
        frame1.data[0]  = 8'h00;  frame1.valid[0]  = 1'b1;  frame1.error[0]  = 1'b0; // Destination Address (01)
        frame1.data[1]  = 8'h00;  frame1.valid[1]  = 1'b1;  frame1.error[1]  = 1'b0;
        frame1.data[2]  = 8'h00;  frame1.valid[2]  = 1'b1;  frame1.error[2]  = 1'b0;
        frame1.data[3]  = 8'h00;  frame1.valid[3]  = 1'b1;  frame1.error[3]  = 1'b0;
        frame1.data[4]  = 8'h00;  frame1.valid[4]  = 1'b1;  frame1.error[4]  = 1'b0;
        frame1.data[5]  = 8'h01;  frame1.valid[5]  = 1'b1;  frame1.error[5]  = 1'b0;
        frame1.data[6]  = 8'h00;  frame1.valid[6]  = 1'b1;  frame1.error[6]  = 1'b0; // Source Address  (02)
        frame1.data[7]  = 8'h00;  frame1.valid[7]  = 1'b1;  frame1.error[7]  = 1'b0;
        frame1.data[8]  = 8'h00;  frame1.valid[8]  = 1'b1;  frame1.error[8]  = 1'b0;
        frame1.data[9]  = 8'h00;  frame1.valid[9]  = 1'b1;  frame1.error[9]  = 1'b0;
        frame1.data[10] = 8'h00;  frame1.valid[10] = 1'b1;  frame1.error[10] = 1'b0;
        frame1.data[11] = 8'h02;  frame1.valid[11] = 1'b1;  frame1.error[11] = 1'b0;
        frame1.data[12] = 8'h81;  frame1.valid[12] = 1'b1;  frame1.error[12] = 1'b0;
        frame1.data[13] = 8'h00;  frame1.valid[13] = 1'b1;  frame1.error[13] = 1'b0; // Length/Type = VLAN

        // VLAN PRI = 7
        frame1.data[  14] = 8'h70; frame1.valid[  14] = 1'b1; frame1.error[  14] = 1'b0;frame1.data[  15] = 8'h00; frame1.valid[  15] = 1'b1; frame1.error[  15] = 1'b0;frame1.data[  16] = 8'h00; frame1.valid[  16] = 1'b1; frame1.error[  16] = 1'b0;frame1.data[  17] = 8'h03; frame1.valid[  17] = 1'b1; frame1.error[  17] = 1'b0;frame1.data[  18] = 8'h04; frame1.valid[  18] = 1'b1; frame1.error[  18] = 1'b0;frame1.data[  19] = 8'h05; frame1.valid[  19] = 1'b1; frame1.error[  19] = 1'b0;frame1.data[  20] = 8'h06; frame1.valid[  20] = 1'b1; frame1.error[  20] = 1'b0;frame1.data[  21] = 8'h07; frame1.valid[  21] = 1'b1; frame1.error[  21] = 1'b0;frame1.data[  22] = 8'h08; frame1.valid[  22] = 1'b1; frame1.error[  22] = 1'b0;frame1.data[  23] = 8'h09; frame1.valid[  23] = 1'b1; frame1.error[  23] = 1'b0;frame1.data[  24] = 8'h0A; frame1.valid[  24] = 1'b1; frame1.error[  24] = 1'b0;frame1.data[  25] = 8'h0B; frame1.valid[  25] = 1'b1; frame1.error[  25] = 1'b0;frame1.data[  26] = 8'h0C; frame1.valid[  26] = 1'b1; frame1.error[  26] = 1'b0;frame1.data[  27] = 8'h0D; frame1.valid[  27] = 1'b1; frame1.error[  27] = 1'b0;frame1.data[  28] = 8'h0E; frame1.valid[  28] = 1'b1; frame1.error[  28] = 1'b0;frame1.data[  29] = 8'h0F; frame1.valid[  29] = 1'b1; frame1.error[  29] = 1'b0;
        frame1.data[  30] = 8'h00; frame1.valid[  30] = 1'b1; frame1.error[  30] = 1'b0;frame1.data[  31] = 8'h11; frame1.valid[  31] = 1'b1; frame1.error[  31] = 1'b0;frame1.data[  32] = 8'h12; frame1.valid[  32] = 1'b1; frame1.error[  32] = 1'b0;frame1.data[  33] = 8'h13; frame1.valid[  33] = 1'b1; frame1.error[  33] = 1'b0;frame1.data[  34] = 8'h00; frame1.valid[  34] = 1'b1; frame1.error[  34] = 1'b0;frame1.data[  35] = 8'h00; frame1.valid[  35] = 1'b1; frame1.error[  35] = 1'b0;frame1.data[  36] = 8'h01; frame1.valid[  36] = 1'b1; frame1.error[  36] = 1'b0;frame1.data[  37] = 8'h02; frame1.valid[  37] = 1'b1; frame1.error[  37] = 1'b0;frame1.data[  38] = 8'h04; frame1.valid[  38] = 1'b1; frame1.error[  38] = 1'b0;frame1.data[  39] = 8'h08; frame1.valid[  39] = 1'b1; frame1.error[  39] = 1'b0;frame1.data[  40] = 8'h10; frame1.valid[  40] = 1'b1; frame1.error[  40] = 1'b0;frame1.data[  41] = 8'h20; frame1.valid[  41] = 1'b1; frame1.error[  41] = 1'b0;frame1.data[  42] = 8'h40; frame1.valid[  42] = 1'b1; frame1.error[  42] = 1'b0;frame1.data[  43] = 8'h80; frame1.valid[  43] = 1'b1; frame1.error[  43] = 1'b0;frame1.data[  44] = 8'h00; frame1.valid[  44] = 1'b1; frame1.error[  44] = 1'b0;frame1.data[  45] = 8'hFF; frame1.valid[  45] = 1'b1; frame1.error[  45] = 1'b0;
        frame1.data[  46] = 8'h10; frame1.valid[  46] = 1'b1; frame1.error[  46] = 1'b0;frame1.data[  47] = 8'h21; frame1.valid[  47] = 1'b1; frame1.error[  47] = 1'b0;frame1.data[  48] = 8'h22; frame1.valid[  48] = 1'b1; frame1.error[  48] = 1'b0;frame1.data[  49] = 8'h23; frame1.valid[  49] = 1'b1; frame1.error[  49] = 1'b0;frame1.data[  50] = 8'h24; frame1.valid[  50] = 1'b1; frame1.error[  50] = 1'b0;frame1.data[  51] = 8'h25; frame1.valid[  51] = 1'b1; frame1.error[  51] = 1'b0;frame1.data[  52] = 8'h26; frame1.valid[  52] = 1'b1; frame1.error[  52] = 1'b0;frame1.data[  53] = 8'h27; frame1.valid[  53] = 1'b1; frame1.error[  53] = 1'b0;frame1.data[  54] = 8'h28; frame1.valid[  54] = 1'b1; frame1.error[  54] = 1'b0;frame1.data[  55] = 8'h29; frame1.valid[  55] = 1'b1; frame1.error[  55] = 1'b0;frame1.data[  56] = 8'h2A; frame1.valid[  56] = 1'b1; frame1.error[  56] = 1'b0;frame1.data[  57] = 8'h2B; frame1.valid[  57] = 1'b1; frame1.error[  57] = 1'b0;frame1.data[  58] = 8'h2C; frame1.valid[  58] = 1'b1; frame1.error[  58] = 1'b0;frame1.data[  59] = 8'h2D; frame1.valid[  59] = 1'b1; frame1.error[  59] = 1'b0;frame1.data[  60] = 8'h2E; frame1.valid[  60] = 1'b1; frame1.error[  60] = 1'b0;frame1.data[  61] = 8'h2F; frame1.valid[  61] = 1'b1; frame1.error[  61] = 1'b0;
        frame1.data[  62] = 8'h00; frame1.valid[  62] = 1'b1; frame1.error[  62] = 1'b0;frame1.data[  63] = 8'h31; frame1.valid[  63] = 1'b1; frame1.error[  63] = 1'b0;frame1.data[  64] = 8'h32; frame1.valid[  64] = 1'b1; frame1.error[  64] = 1'b0;frame1.data[  65] = 8'h33; frame1.valid[  65] = 1'b1; frame1.error[  65] = 1'b0;frame1.data[  66] = 8'h34; frame1.valid[  66] = 1'b1; frame1.error[  66] = 1'b0;frame1.data[  67] = 8'h35; frame1.valid[  67] = 1'b1; frame1.error[  67] = 1'b0;frame1.data[  68] = 8'h36; frame1.valid[  68] = 1'b1; frame1.error[  68] = 1'b0;frame1.data[  69] = 8'h37; frame1.valid[  69] = 1'b1; frame1.error[  69] = 1'b0;frame1.data[  70] = 8'h38; frame1.valid[  70] = 1'b1; frame1.error[  70] = 1'b0;frame1.data[  71] = 8'h39; frame1.valid[  71] = 1'b1; frame1.error[  71] = 1'b0;frame1.data[  72] = 8'h3A; frame1.valid[  72] = 1'b1; frame1.error[  72] = 1'b0;frame1.data[  73] = 8'h3B; frame1.valid[  73] = 1'b1; frame1.error[  73] = 1'b0;frame1.data[  74] = 8'h3C; frame1.valid[  74] = 1'b1; frame1.error[  74] = 1'b0;frame1.data[  75] = 8'h3D; frame1.valid[  75] = 1'b1; frame1.error[  75] = 1'b0;frame1.data[  76] = 8'h3E; frame1.valid[  76] = 1'b1; frame1.error[  76] = 1'b0;frame1.data[  77] = 8'h3F; frame1.valid[  77] = 1'b1; frame1.error[  77] = 1'b0;
        frame1.data[  78] = 8'h00; frame1.valid[  78] = 1'b1; frame1.error[  78] = 1'b0;frame1.data[  79] = 8'h41; frame1.valid[  79] = 1'b1; frame1.error[  79] = 1'b0;frame1.data[  80] = 8'h42; frame1.valid[  80] = 1'b1; frame1.error[  80] = 1'b0;frame1.data[  81] = 8'h43; frame1.valid[  81] = 1'b1; frame1.error[  81] = 1'b0;frame1.data[  82] = 8'h44; frame1.valid[  82] = 1'b1; frame1.error[  82] = 1'b0;frame1.data[  83] = 8'h45; frame1.valid[  83] = 1'b1; frame1.error[  83] = 1'b0;frame1.data[  84] = 8'h46; frame1.valid[  84] = 1'b1; frame1.error[  84] = 1'b0;frame1.data[  85] = 8'h47; frame1.valid[  85] = 1'b1; frame1.error[  85] = 1'b0;frame1.data[  86] = 8'h48; frame1.valid[  86] = 1'b1; frame1.error[  86] = 1'b0;frame1.data[  87] = 8'h49; frame1.valid[  87] = 1'b1; frame1.error[  87] = 1'b0;frame1.data[  88] = 8'h4A; frame1.valid[  88] = 1'b1; frame1.error[  88] = 1'b0;frame1.data[  89] = 8'h4B; frame1.valid[  89] = 1'b1; frame1.error[  89] = 1'b0;frame1.data[  90] = 8'h4C; frame1.valid[  90] = 1'b1; frame1.error[  90] = 1'b0;frame1.data[  91] = 8'h4D; frame1.valid[  91] = 1'b1; frame1.error[  91] = 1'b0;frame1.data[  92] = 8'h4E; frame1.valid[  92] = 1'b1; frame1.error[  92] = 1'b0;frame1.data[  93] = 8'h4F; frame1.valid[  93] = 1'b1; frame1.error[  93] = 1'b0;
        frame1.data[  94] = 8'h00; frame1.valid[  94] = 1'b1; frame1.error[  94] = 1'b0;frame1.data[  95] = 8'h51; frame1.valid[  95] = 1'b1; frame1.error[  95] = 1'b0;frame1.data[  96] = 8'h52; frame1.valid[  96] = 1'b1; frame1.error[  96] = 1'b0;frame1.data[  97] = 8'h53; frame1.valid[  97] = 1'b1; frame1.error[  97] = 1'b0;frame1.data[  98] = 8'h54; frame1.valid[  98] = 1'b1; frame1.error[  98] = 1'b0;frame1.data[  99] = 8'h55; frame1.valid[  99] = 1'b1; frame1.error[  99] = 1'b0;frame1.data[ 100] = 8'h56; frame1.valid[ 100] = 1'b1; frame1.error[ 100] = 1'b0;frame1.data[ 101] = 8'h57; frame1.valid[ 101] = 1'b1; frame1.error[ 101] = 1'b0;frame1.data[ 102] = 8'h58; frame1.valid[ 102] = 1'b1; frame1.error[ 102] = 1'b0;frame1.data[ 103] = 8'h59; frame1.valid[ 103] = 1'b1; frame1.error[ 103] = 1'b0;frame1.data[ 104] = 8'h5A; frame1.valid[ 104] = 1'b1; frame1.error[ 104] = 1'b0;frame1.data[ 105] = 8'h5B; frame1.valid[ 105] = 1'b1; frame1.error[ 105] = 1'b0;frame1.data[ 106] = 8'h5C; frame1.valid[ 106] = 1'b1; frame1.error[ 106] = 1'b0;frame1.data[ 107] = 8'h5D; frame1.valid[ 107] = 1'b1; frame1.error[ 107] = 1'b0;frame1.data[ 108] = 8'h5E; frame1.valid[ 108] = 1'b1; frame1.error[ 108] = 1'b0;frame1.data[ 109] = 8'h5F; frame1.valid[ 109] = 1'b1; frame1.error[ 109] = 1'b0;
        frame1.data[ 110] = 8'h00; frame1.valid[ 110] = 1'b1; frame1.error[ 110] = 1'b0;frame1.data[ 111] = 8'h61; frame1.valid[ 111] = 1'b1; frame1.error[ 111] = 1'b0;frame1.data[ 112] = 8'h62; frame1.valid[ 112] = 1'b1; frame1.error[ 112] = 1'b0;frame1.data[ 113] = 8'h63; frame1.valid[ 113] = 1'b1; frame1.error[ 113] = 1'b0;frame1.data[ 114] = 8'h64; frame1.valid[ 114] = 1'b1; frame1.error[ 114] = 1'b0;frame1.data[ 115] = 8'h65; frame1.valid[ 115] = 1'b1; frame1.error[ 115] = 1'b0;frame1.data[ 116] = 8'h66; frame1.valid[ 116] = 1'b1; frame1.error[ 116] = 1'b0;frame1.data[ 117] = 8'h67; frame1.valid[ 117] = 1'b1; frame1.error[ 117] = 1'b0;frame1.data[ 118] = 8'h68; frame1.valid[ 118] = 1'b1; frame1.error[ 118] = 1'b0;frame1.data[ 119] = 8'h69; frame1.valid[ 119] = 1'b1; frame1.error[ 119] = 1'b0;frame1.data[ 120] = 8'h6A; frame1.valid[ 120] = 1'b1; frame1.error[ 120] = 1'b0;frame1.data[ 121] = 8'h6B; frame1.valid[ 121] = 1'b1; frame1.error[ 121] = 1'b0;frame1.data[ 122] = 8'h6C; frame1.valid[ 122] = 1'b1; frame1.error[ 122] = 1'b0;frame1.data[ 123] = 8'h6D; frame1.valid[ 123] = 1'b1; frame1.error[ 123] = 1'b0;frame1.data[ 124] = 8'h6E; frame1.valid[ 124] = 1'b1; frame1.error[ 124] = 1'b0;frame1.data[ 125] = 8'h6F; frame1.valid[ 125] = 1'b1; frame1.error[ 125] = 1'b0;
        frame1.data[ 126] = 8'h00; frame1.valid[ 126] = 1'b1; frame1.error[ 126] = 1'b0;frame1.data[ 127] = 8'h71; frame1.valid[ 127] = 1'b1; frame1.error[ 127] = 1'b0;frame1.data[ 128] = 8'h72; frame1.valid[ 128] = 1'b1; frame1.error[ 128] = 1'b0;frame1.data[ 129] = 8'h73; frame1.valid[ 129] = 1'b1; frame1.error[ 129] = 1'b0;frame1.data[ 130] = 8'h74; frame1.valid[ 130] = 1'b1; frame1.error[ 130] = 1'b0;frame1.data[ 131] = 8'h75; frame1.valid[ 131] = 1'b1; frame1.error[ 131] = 1'b0;frame1.data[ 132] = 8'h76; frame1.valid[ 132] = 1'b1; frame1.error[ 132] = 1'b0;frame1.data[ 133] = 8'h77; frame1.valid[ 133] = 1'b1; frame1.error[ 133] = 1'b0;frame1.data[ 134] = 8'h78; frame1.valid[ 134] = 1'b1; frame1.error[ 134] = 1'b0;frame1.data[ 135] = 8'h79; frame1.valid[ 135] = 1'b1; frame1.error[ 135] = 1'b0;frame1.data[ 136] = 8'h7A; frame1.valid[ 136] = 1'b1; frame1.error[ 136] = 1'b0;frame1.data[ 137] = 8'h7B; frame1.valid[ 137] = 1'b1; frame1.error[ 137] = 1'b0;frame1.data[ 138] = 8'h7C; frame1.valid[ 138] = 1'b1; frame1.error[ 138] = 1'b0;frame1.data[ 139] = 8'h7D; frame1.valid[ 139] = 1'b1; frame1.error[ 139] = 1'b0;frame1.data[ 140] = 8'h7E; frame1.valid[ 140] = 1'b1; frame1.error[ 140] = 1'b0;frame1.data[ 141] = 8'h7F; frame1.valid[ 141] = 1'b1; frame1.error[ 141] = 1'b0;
        frame1.data[ 142] = 8'h00; frame1.valid[ 142] = 1'b1; frame1.error[ 142] = 1'b0;frame1.data[ 143] = 8'h81; frame1.valid[ 143] = 1'b1; frame1.error[ 143] = 1'b0;frame1.data[ 144] = 8'h82; frame1.valid[ 144] = 1'b1; frame1.error[ 144] = 1'b0;frame1.data[ 145] = 8'h83; frame1.valid[ 145] = 1'b1; frame1.error[ 145] = 1'b0;frame1.data[ 146] = 8'h84; frame1.valid[ 146] = 1'b1; frame1.error[ 146] = 1'b0;frame1.data[ 147] = 8'h85; frame1.valid[ 147] = 1'b1; frame1.error[ 147] = 1'b0;frame1.data[ 148] = 8'h86; frame1.valid[ 148] = 1'b1; frame1.error[ 148] = 1'b0;frame1.data[ 149] = 8'h87; frame1.valid[ 149] = 1'b1; frame1.error[ 149] = 1'b0;frame1.data[ 150] = 8'h88; frame1.valid[ 150] = 1'b1; frame1.error[ 150] = 1'b0;frame1.data[ 151] = 8'h89; frame1.valid[ 151] = 1'b1; frame1.error[ 151] = 1'b0;frame1.data[ 152] = 8'h8A; frame1.valid[ 152] = 1'b1; frame1.error[ 152] = 1'b0;frame1.data[ 153] = 8'h8B; frame1.valid[ 153] = 1'b1; frame1.error[ 153] = 1'b0;frame1.data[ 154] = 8'h8C; frame1.valid[ 154] = 1'b1; frame1.error[ 154] = 1'b0;frame1.data[ 155] = 8'h8D; frame1.valid[ 155] = 1'b1; frame1.error[ 155] = 1'b0;frame1.data[ 156] = 8'h8E; frame1.valid[ 156] = 1'b1; frame1.error[ 156] = 1'b0;frame1.data[ 157] = 8'h8F; frame1.valid[ 157] = 1'b1; frame1.error[ 157] = 1'b0;
        frame1.data[ 158] = 8'h00; frame1.valid[ 158] = 1'b1; frame1.error[ 158] = 1'b0;frame1.data[ 159] = 8'h91; frame1.valid[ 159] = 1'b1; frame1.error[ 159] = 1'b0;frame1.data[ 160] = 8'h92; frame1.valid[ 160] = 1'b1; frame1.error[ 160] = 1'b0;frame1.data[ 161] = 8'h93; frame1.valid[ 161] = 1'b1; frame1.error[ 161] = 1'b0;frame1.data[ 162] = 8'h94; frame1.valid[ 162] = 1'b1; frame1.error[ 162] = 1'b0;frame1.data[ 163] = 8'h95; frame1.valid[ 163] = 1'b1; frame1.error[ 163] = 1'b0;frame1.data[ 164] = 8'h96; frame1.valid[ 164] = 1'b1; frame1.error[ 164] = 1'b0;frame1.data[ 165] = 8'h97; frame1.valid[ 165] = 1'b1; frame1.error[ 165] = 1'b0;frame1.data[ 166] = 8'h98; frame1.valid[ 166] = 1'b1; frame1.error[ 166] = 1'b0;frame1.data[ 167] = 8'h99; frame1.valid[ 167] = 1'b1; frame1.error[ 167] = 1'b0;frame1.data[ 168] = 8'h9A; frame1.valid[ 168] = 1'b1; frame1.error[ 168] = 1'b0;frame1.data[ 169] = 8'h9B; frame1.valid[ 169] = 1'b1; frame1.error[ 169] = 1'b0;frame1.data[ 170] = 8'h9C; frame1.valid[ 170] = 1'b1; frame1.error[ 170] = 1'b0;frame1.data[ 171] = 8'h9D; frame1.valid[ 171] = 1'b1; frame1.error[ 171] = 1'b0;frame1.data[ 172] = 8'h9E; frame1.valid[ 172] = 1'b1; frame1.error[ 172] = 1'b0;frame1.data[ 173] = 8'h9F; frame1.valid[ 173] = 1'b1; frame1.error[ 173] = 1'b0;
        frame1.data[ 174] = 8'hA0; frame1.valid[ 174] = 1'b1; frame1.error[ 174] = 1'b0;frame1.data[ 175] = 8'hA1; frame1.valid[ 175] = 1'b1; frame1.error[ 175] = 1'b0;frame1.data[ 176] = 8'hA2; frame1.valid[ 176] = 1'b1; frame1.error[ 176] = 1'b0;frame1.data[ 177] = 8'hA3; frame1.valid[ 177] = 1'b1; frame1.error[ 177] = 1'b0;frame1.data[ 178] = 8'hA4; frame1.valid[ 178] = 1'b1; frame1.error[ 178] = 1'b0;frame1.data[ 179] = 8'hA5; frame1.valid[ 179] = 1'b1; frame1.error[ 179] = 1'b0;frame1.data[ 180] = 8'hA6; frame1.valid[ 180] = 1'b1; frame1.error[ 180] = 1'b0;frame1.data[ 181] = 8'hA7; frame1.valid[ 181] = 1'b1; frame1.error[ 181] = 1'b0;frame1.data[ 182] = 8'hA8; frame1.valid[ 182] = 1'b1; frame1.error[ 182] = 1'b0;frame1.data[ 183] = 8'hA9; frame1.valid[ 183] = 1'b1; frame1.error[ 183] = 1'b0;frame1.data[ 184] = 8'hAA; frame1.valid[ 184] = 1'b1; frame1.error[ 184] = 1'b0;frame1.data[ 185] = 8'hAB; frame1.valid[ 185] = 1'b1; frame1.error[ 185] = 1'b0;frame1.data[ 186] = 8'hAC; frame1.valid[ 186] = 1'b1; frame1.error[ 186] = 1'b0;frame1.data[ 187] = 8'hAD; frame1.valid[ 187] = 1'b1; frame1.error[ 187] = 1'b0;frame1.data[ 188] = 8'hAE; frame1.valid[ 188] = 1'b1; frame1.error[ 188] = 1'b0;frame1.data[ 189] = 8'hAF; frame1.valid[ 189] = 1'b1; frame1.error[ 189] = 1'b0;
        frame1.data[ 190] = 8'hB0; frame1.valid[ 190] = 1'b1; frame1.error[ 190] = 1'b0;frame1.data[ 191] = 8'hB1; frame1.valid[ 191] = 1'b1; frame1.error[ 191] = 1'b0;frame1.data[ 192] = 8'hB2; frame1.valid[ 192] = 1'b1; frame1.error[ 192] = 1'b0;frame1.data[ 193] = 8'hB3; frame1.valid[ 193] = 1'b1; frame1.error[ 193] = 1'b0;frame1.data[ 194] = 8'hB4; frame1.valid[ 194] = 1'b1; frame1.error[ 194] = 1'b0;frame1.data[ 195] = 8'hB5; frame1.valid[ 195] = 1'b1; frame1.error[ 195] = 1'b0;frame1.data[ 196] = 8'hB6; frame1.valid[ 196] = 1'b1; frame1.error[ 196] = 1'b0;frame1.data[ 197] = 8'hB7; frame1.valid[ 197] = 1'b1; frame1.error[ 197] = 1'b0;frame1.data[ 198] = 8'hB8; frame1.valid[ 198] = 1'b1; frame1.error[ 198] = 1'b0;frame1.data[ 199] = 8'hB9; frame1.valid[ 199] = 1'b1; frame1.error[ 199] = 1'b0;frame1.data[ 200] = 8'hBA; frame1.valid[ 200] = 1'b1; frame1.error[ 200] = 1'b0;frame1.data[ 201] = 8'hBB; frame1.valid[ 201] = 1'b1; frame1.error[ 201] = 1'b0;frame1.data[ 202] = 8'hBC; frame1.valid[ 202] = 1'b1; frame1.error[ 202] = 1'b0;frame1.data[ 203] = 8'hBD; frame1.valid[ 203] = 1'b1; frame1.error[ 203] = 1'b0;frame1.data[ 204] = 8'hBE; frame1.valid[ 204] = 1'b1; frame1.error[ 204] = 1'b0;frame1.data[ 205] = 8'hBF; frame1.valid[ 205] = 1'b1; frame1.error[ 205] = 1'b0;
        frame1.data[ 206] = 8'hC0; frame1.valid[ 206] = 1'b1; frame1.error[ 206] = 1'b0;frame1.data[ 207] = 8'hC1; frame1.valid[ 207] = 1'b1; frame1.error[ 207] = 1'b0;frame1.data[ 208] = 8'hC2; frame1.valid[ 208] = 1'b1; frame1.error[ 208] = 1'b0;frame1.data[ 209] = 8'hC3; frame1.valid[ 209] = 1'b1; frame1.error[ 209] = 1'b0;frame1.data[ 210] = 8'hC4; frame1.valid[ 210] = 1'b1; frame1.error[ 210] = 1'b0;frame1.data[ 211] = 8'hC5; frame1.valid[ 211] = 1'b1; frame1.error[ 211] = 1'b0;frame1.data[ 212] = 8'hC6; frame1.valid[ 212] = 1'b1; frame1.error[ 212] = 1'b0;frame1.data[ 213] = 8'hC7; frame1.valid[ 213] = 1'b1; frame1.error[ 213] = 1'b0;frame1.data[ 214] = 8'hC8; frame1.valid[ 214] = 1'b1; frame1.error[ 214] = 1'b0;frame1.data[ 215] = 8'hC9; frame1.valid[ 215] = 1'b1; frame1.error[ 215] = 1'b0;frame1.data[ 216] = 8'hCA; frame1.valid[ 216] = 1'b1; frame1.error[ 216] = 1'b0;frame1.data[ 217] = 8'hCB; frame1.valid[ 217] = 1'b1; frame1.error[ 217] = 1'b0;frame1.data[ 218] = 8'hCC; frame1.valid[ 218] = 1'b1; frame1.error[ 218] = 1'b0;frame1.data[ 219] = 8'hCD; frame1.valid[ 219] = 1'b1; frame1.error[ 219] = 1'b0;frame1.data[ 220] = 8'hCE; frame1.valid[ 220] = 1'b1; frame1.error[ 220] = 1'b0;frame1.data[ 221] = 8'hCF; frame1.valid[ 221] = 1'b1; frame1.error[ 221] = 1'b0;
        frame1.data[ 222] = 8'hD0; frame1.valid[ 222] = 1'b1; frame1.error[ 222] = 1'b0;frame1.data[ 223] = 8'hD1; frame1.valid[ 223] = 1'b1; frame1.error[ 223] = 1'b0;frame1.data[ 224] = 8'hD2; frame1.valid[ 224] = 1'b1; frame1.error[ 224] = 1'b0;frame1.data[ 225] = 8'hD3; frame1.valid[ 225] = 1'b1; frame1.error[ 225] = 1'b0;frame1.data[ 226] = 8'hD4; frame1.valid[ 226] = 1'b1; frame1.error[ 226] = 1'b0;frame1.data[ 227] = 8'hD5; frame1.valid[ 227] = 1'b1; frame1.error[ 227] = 1'b0;frame1.data[ 228] = 8'hD6; frame1.valid[ 228] = 1'b1; frame1.error[ 228] = 1'b0;frame1.data[ 229] = 8'hD7; frame1.valid[ 229] = 1'b1; frame1.error[ 229] = 1'b0;frame1.data[ 230] = 8'hD8; frame1.valid[ 230] = 1'b1; frame1.error[ 230] = 1'b0;frame1.data[ 231] = 8'hD9; frame1.valid[ 231] = 1'b1; frame1.error[ 231] = 1'b0;frame1.data[ 232] = 8'hDA; frame1.valid[ 232] = 1'b1; frame1.error[ 232] = 1'b0;frame1.data[ 233] = 8'hDB; frame1.valid[ 233] = 1'b1; frame1.error[ 233] = 1'b0;frame1.data[ 234] = 8'hDC; frame1.valid[ 234] = 1'b1; frame1.error[ 234] = 1'b0;frame1.data[ 235] = 8'hDD; frame1.valid[ 235] = 1'b1; frame1.error[ 235] = 1'b0;frame1.data[ 236] = 8'hDE; frame1.valid[ 236] = 1'b1; frame1.error[ 236] = 1'b0;frame1.data[ 237] = 8'hDF; frame1.valid[ 237] = 1'b1; frame1.error[ 237] = 1'b0;
        frame1.data[ 238] = 8'hE0; frame1.valid[ 238] = 1'b1; frame1.error[ 238] = 1'b0;frame1.data[ 239] = 8'hE1; frame1.valid[ 239] = 1'b1; frame1.error[ 239] = 1'b0;frame1.data[ 240] = 8'hE2; frame1.valid[ 240] = 1'b1; frame1.error[ 240] = 1'b0;frame1.data[ 241] = 8'hE3; frame1.valid[ 241] = 1'b1; frame1.error[ 241] = 1'b0;frame1.data[ 242] = 8'hE4; frame1.valid[ 242] = 1'b1; frame1.error[ 242] = 1'b0;frame1.data[ 243] = 8'hE5; frame1.valid[ 243] = 1'b1; frame1.error[ 243] = 1'b0;frame1.data[ 244] = 8'hE6; frame1.valid[ 244] = 1'b1; frame1.error[ 244] = 1'b0;frame1.data[ 245] = 8'hE7; frame1.valid[ 245] = 1'b1; frame1.error[ 245] = 1'b0;frame1.data[ 246] = 8'hE8; frame1.valid[ 246] = 1'b1; frame1.error[ 246] = 1'b0;frame1.data[ 247] = 8'hE9; frame1.valid[ 247] = 1'b1; frame1.error[ 247] = 1'b0;frame1.data[ 248] = 8'hEA; frame1.valid[ 248] = 1'b1; frame1.error[ 248] = 1'b0;frame1.data[ 249] = 8'hEB; frame1.valid[ 249] = 1'b1; frame1.error[ 249] = 1'b0;frame1.data[ 250] = 8'hEC; frame1.valid[ 250] = 1'b1; frame1.error[ 250] = 1'b0;frame1.data[ 251] = 8'hED; frame1.valid[ 251] = 1'b1; frame1.error[ 251] = 1'b0;frame1.data[ 252] = 8'hEE; frame1.valid[ 252] = 1'b1; frame1.error[ 252] = 1'b0;frame1.data[ 253] = 8'hEF; frame1.valid[ 253] = 1'b1; frame1.error[ 253] = 1'b0;
        frame1.data[ 254] = 8'hF0; frame1.valid[ 254] = 1'b1; frame1.error[ 254] = 1'b0;frame1.data[ 255] = 8'hF1; frame1.valid[ 255] = 1'b1; frame1.error[ 255] = 1'b0;frame1.data[ 256] = 8'hF2; frame1.valid[ 256] = 1'b1; frame1.error[ 256] = 1'b0;frame1.data[ 257] = 8'hF3; frame1.valid[ 257] = 1'b1; frame1.error[ 257] = 1'b0;frame1.data[ 258] = 8'hF4; frame1.valid[ 258] = 1'b1; frame1.error[ 258] = 1'b0;frame1.data[ 259] = 8'hF5; frame1.valid[ 259] = 1'b1; frame1.error[ 259] = 1'b0;frame1.data[ 260] = 8'hF6; frame1.valid[ 260] = 1'b1; frame1.error[ 260] = 1'b0;frame1.data[ 261] = 8'hF7; frame1.valid[ 261] = 1'b1; frame1.error[ 261] = 1'b0;frame1.data[ 262] = 8'hF8; frame1.valid[ 262] = 1'b1; frame1.error[ 262] = 1'b0;frame1.data[ 263] = 8'hF9; frame1.valid[ 263] = 1'b1; frame1.error[ 263] = 1'b0;frame1.data[ 264] = 8'hFA; frame1.valid[ 264] = 1'b1; frame1.error[ 264] = 1'b0;frame1.data[ 265] = 8'hFB; frame1.valid[ 265] = 1'b1; frame1.error[ 265] = 1'b0;frame1.data[ 266] = 8'hFC; frame1.valid[ 266] = 1'b1; frame1.error[ 266] = 1'b0;frame1.data[ 267] = 8'hFD; frame1.valid[ 267] = 1'b1; frame1.error[ 267] = 1'b0;frame1.data[ 268] = 8'hFE; frame1.valid[ 268] = 1'b1; frame1.error[ 268] = 1'b0;frame1.data[ 269] = 8'h00; frame1.valid[ 269] = 1'b1; frame1.error[ 269] = 1'b0;
        frame1.data[ 270] = 8'h01; frame1.valid[ 270] = 1'b1; frame1.error[ 270] = 1'b0;frame1.data[ 271] = 8'h02; frame1.valid[ 271] = 1'b1; frame1.error[ 271] = 1'b0;frame1.data[ 272] = 8'h03; frame1.valid[ 272] = 1'b1; frame1.error[ 272] = 1'b0;frame1.data[ 273] = 8'h04; frame1.valid[ 273] = 1'b1; frame1.error[ 273] = 1'b0;frame1.data[ 274] = 8'h05; frame1.valid[ 274] = 1'b1; frame1.error[ 274] = 1'b0;frame1.data[ 275] = 8'h06; frame1.valid[ 275] = 1'b1; frame1.error[ 275] = 1'b0;frame1.data[ 276] = 8'h07; frame1.valid[ 276] = 1'b1; frame1.error[ 276] = 1'b0;frame1.data[ 277] = 8'h08; frame1.valid[ 277] = 1'b1; frame1.error[ 277] = 1'b0;frame1.data[ 278] = 8'h09; frame1.valid[ 278] = 1'b1; frame1.error[ 278] = 1'b0;frame1.data[ 279] = 8'h0A; frame1.valid[ 279] = 1'b1; frame1.error[ 279] = 1'b0;frame1.data[ 280] = 8'h0B; frame1.valid[ 280] = 1'b1; frame1.error[ 280] = 1'b0;frame1.data[ 281] = 8'h0C; frame1.valid[ 281] = 1'b1; frame1.error[ 281] = 1'b0;frame1.data[ 282] = 8'h0D; frame1.valid[ 282] = 1'b1; frame1.error[ 282] = 1'b0;frame1.data[ 283] = 8'h0E; frame1.valid[ 283] = 1'b1; frame1.error[ 283] = 1'b0;frame1.data[ 284] = 8'h0F; frame1.valid[ 284] = 1'b1; frame1.error[ 284] = 1'b0;frame1.data[ 285] = 8'h10; frame1.valid[ 285] = 1'b1; frame1.error[ 285] = 1'b0;
        frame1.data[ 286] = 8'h11; frame1.valid[ 286] = 1'b1; frame1.error[ 286] = 1'b0;frame1.data[ 287] = 8'h12; frame1.valid[ 287] = 1'b1; frame1.error[ 287] = 1'b0;frame1.data[ 288] = 8'h13; frame1.valid[ 288] = 1'b1; frame1.error[ 288] = 1'b0;frame1.data[ 289] = 8'h14; frame1.valid[ 289] = 1'b1; frame1.error[ 289] = 1'b0;frame1.data[ 290] = 8'h15; frame1.valid[ 290] = 1'b1; frame1.error[ 290] = 1'b0;frame1.data[ 291] = 8'h16; frame1.valid[ 291] = 1'b1; frame1.error[ 291] = 1'b0;frame1.data[ 292] = 8'h17; frame1.valid[ 292] = 1'b1; frame1.error[ 292] = 1'b0;frame1.data[ 293] = 8'h18; frame1.valid[ 293] = 1'b1; frame1.error[ 293] = 1'b0;frame1.data[ 294] = 8'h19; frame1.valid[ 294] = 1'b1; frame1.error[ 294] = 1'b0;frame1.data[ 295] = 8'h1A; frame1.valid[ 295] = 1'b1; frame1.error[ 295] = 1'b0;frame1.data[ 296] = 8'h1B; frame1.valid[ 296] = 1'b1; frame1.error[ 296] = 1'b0;frame1.data[ 297] = 8'h1C; frame1.valid[ 297] = 1'b1; frame1.error[ 297] = 1'b0;frame1.data[ 298] = 8'h1D; frame1.valid[ 298] = 1'b1; frame1.error[ 298] = 1'b0;frame1.data[ 299] = 8'h1E; frame1.valid[ 299] = 1'b1; frame1.error[ 299] = 1'b0;frame1.data[ 300] = 8'h1F; frame1.valid[ 300] = 1'b1; frame1.error[ 300] = 1'b0;frame1.data[ 301] = 8'h20; frame1.valid[ 301] = 1'b1; frame1.error[ 301] = 1'b0;
        frame1.data[ 302] = 8'h21; frame1.valid[ 302] = 1'b1; frame1.error[ 302] = 1'b0;frame1.data[ 303] = 8'h22; frame1.valid[ 303] = 1'b1; frame1.error[ 303] = 1'b0;frame1.data[ 304] = 8'h23; frame1.valid[ 304] = 1'b1; frame1.error[ 304] = 1'b0;frame1.data[ 305] = 8'h24; frame1.valid[ 305] = 1'b1; frame1.error[ 305] = 1'b0;frame1.data[ 306] = 8'h25; frame1.valid[ 306] = 1'b1; frame1.error[ 306] = 1'b0;frame1.data[ 307] = 8'h26; frame1.valid[ 307] = 1'b1; frame1.error[ 307] = 1'b0;frame1.data[ 308] = 8'h27; frame1.valid[ 308] = 1'b1; frame1.error[ 308] = 1'b0;frame1.data[ 309] = 8'h28; frame1.valid[ 309] = 1'b1; frame1.error[ 309] = 1'b0;frame1.data[ 310] = 8'h29; frame1.valid[ 310] = 1'b1; frame1.error[ 310] = 1'b0;frame1.data[ 311] = 8'h2A; frame1.valid[ 311] = 1'b1; frame1.error[ 311] = 1'b0;frame1.data[ 312] = 8'h2B; frame1.valid[ 312] = 1'b1; frame1.error[ 312] = 1'b0;frame1.data[ 313] = 8'h2C; frame1.valid[ 313] = 1'b1; frame1.error[ 313] = 1'b0;frame1.data[ 314] = 8'h2D; frame1.valid[ 314] = 1'b1; frame1.error[ 314] = 1'b0;frame1.data[ 315] = 8'h2E; frame1.valid[ 315] = 1'b1; frame1.error[ 315] = 1'b0;frame1.data[ 316] = 8'h2F; frame1.valid[ 316] = 1'b1; frame1.error[ 316] = 1'b0;frame1.data[ 317] = 8'h30; frame1.valid[ 317] = 1'b1; frame1.error[ 317] = 1'b0;
        frame1.data[ 318] = 8'h31; frame1.valid[ 318] = 1'b1; frame1.error[ 318] = 1'b0;frame1.data[ 319] = 8'h32; frame1.valid[ 319] = 1'b1; frame1.error[ 319] = 1'b0;frame1.data[ 320] = 8'h33; frame1.valid[ 320] = 1'b1; frame1.error[ 320] = 1'b0;frame1.data[ 321] = 8'h34; frame1.valid[ 321] = 1'b1; frame1.error[ 321] = 1'b0;frame1.data[ 322] = 8'h35; frame1.valid[ 322] = 1'b1; frame1.error[ 322] = 1'b0;frame1.data[ 323] = 8'h36; frame1.valid[ 323] = 1'b1; frame1.error[ 323] = 1'b0;frame1.data[ 324] = 8'h37; frame1.valid[ 324] = 1'b1; frame1.error[ 324] = 1'b0;frame1.data[ 325] = 8'h38; frame1.valid[ 325] = 1'b1; frame1.error[ 325] = 1'b0;frame1.data[ 326] = 8'h39; frame1.valid[ 326] = 1'b1; frame1.error[ 326] = 1'b0;frame1.data[ 327] = 8'h3A; frame1.valid[ 327] = 1'b1; frame1.error[ 327] = 1'b0;frame1.data[ 328] = 8'h3B; frame1.valid[ 328] = 1'b1; frame1.error[ 328] = 1'b0;frame1.data[ 329] = 8'h3C; frame1.valid[ 329] = 1'b1; frame1.error[ 329] = 1'b0;frame1.data[ 330] = 8'h3D; frame1.valid[ 330] = 1'b1; frame1.error[ 330] = 1'b0;frame1.data[ 331] = 8'h3E; frame1.valid[ 331] = 1'b1; frame1.error[ 331] = 1'b0;frame1.data[ 332] = 8'h3F; frame1.valid[ 332] = 1'b1; frame1.error[ 332] = 1'b0;frame1.data[ 333] = 8'h40; frame1.valid[ 333] = 1'b1; frame1.error[ 333] = 1'b0;
        frame1.data[ 334] = 8'h41; frame1.valid[ 334] = 1'b1; frame1.error[ 334] = 1'b0;frame1.data[ 335] = 8'h42; frame1.valid[ 335] = 1'b1; frame1.error[ 335] = 1'b0;frame1.data[ 336] = 8'h43; frame1.valid[ 336] = 1'b1; frame1.error[ 336] = 1'b0;frame1.data[ 337] = 8'h44; frame1.valid[ 337] = 1'b1; frame1.error[ 337] = 1'b0;frame1.data[ 338] = 8'h45; frame1.valid[ 338] = 1'b1; frame1.error[ 338] = 1'b0;frame1.data[ 339] = 8'h46; frame1.valid[ 339] = 1'b1; frame1.error[ 339] = 1'b0;frame1.data[ 340] = 8'h47; frame1.valid[ 340] = 1'b1; frame1.error[ 340] = 1'b0;frame1.data[ 341] = 8'h48; frame1.valid[ 341] = 1'b1; frame1.error[ 341] = 1'b0;frame1.data[ 342] = 8'h49; frame1.valid[ 342] = 1'b1; frame1.error[ 342] = 1'b0;frame1.data[ 343] = 8'h4A; frame1.valid[ 343] = 1'b1; frame1.error[ 343] = 1'b0;frame1.data[ 344] = 8'h4B; frame1.valid[ 344] = 1'b1; frame1.error[ 344] = 1'b0;frame1.data[ 345] = 8'h4C; frame1.valid[ 345] = 1'b1; frame1.error[ 345] = 1'b0;frame1.data[ 346] = 8'h4D; frame1.valid[ 346] = 1'b1; frame1.error[ 346] = 1'b0;frame1.data[ 347] = 8'h4E; frame1.valid[ 347] = 1'b1; frame1.error[ 347] = 1'b0;frame1.data[ 348] = 8'h4F; frame1.valid[ 348] = 1'b1; frame1.error[ 348] = 1'b0;frame1.data[ 349] = 8'h50; frame1.valid[ 349] = 1'b1; frame1.error[ 349] = 1'b0;
        frame1.data[ 350] = 8'h51; frame1.valid[ 350] = 1'b1; frame1.error[ 350] = 1'b0;frame1.data[ 351] = 8'h52; frame1.valid[ 351] = 1'b1; frame1.error[ 351] = 1'b0;frame1.data[ 352] = 8'h53; frame1.valid[ 352] = 1'b1; frame1.error[ 352] = 1'b0;frame1.data[ 353] = 8'h54; frame1.valid[ 353] = 1'b1; frame1.error[ 353] = 1'b0;frame1.data[ 354] = 8'h55; frame1.valid[ 354] = 1'b1; frame1.error[ 354] = 1'b0;frame1.data[ 355] = 8'h56; frame1.valid[ 355] = 1'b1; frame1.error[ 355] = 1'b0;frame1.data[ 356] = 8'h57; frame1.valid[ 356] = 1'b1; frame1.error[ 356] = 1'b0;frame1.data[ 357] = 8'h58; frame1.valid[ 357] = 1'b1; frame1.error[ 357] = 1'b0;frame1.data[ 358] = 8'h59; frame1.valid[ 358] = 1'b1; frame1.error[ 358] = 1'b0;frame1.data[ 359] = 8'h5A; frame1.valid[ 359] = 1'b1; frame1.error[ 359] = 1'b0;frame1.data[ 360] = 8'h5B; frame1.valid[ 360] = 1'b1; frame1.error[ 360] = 1'b0;frame1.data[ 361] = 8'h5C; frame1.valid[ 361] = 1'b1; frame1.error[ 361] = 1'b0;frame1.data[ 362] = 8'h5D; frame1.valid[ 362] = 1'b1; frame1.error[ 362] = 1'b0;frame1.data[ 363] = 8'h5E; frame1.valid[ 363] = 1'b1; frame1.error[ 363] = 1'b0;frame1.data[ 364] = 8'h5F; frame1.valid[ 364] = 1'b1; frame1.error[ 364] = 1'b0;frame1.data[ 365] = 8'h60; frame1.valid[ 365] = 1'b1; frame1.error[ 365] = 1'b0;
        frame1.data[ 366] = 8'h61; frame1.valid[ 366] = 1'b1; frame1.error[ 366] = 1'b0;frame1.data[ 367] = 8'h62; frame1.valid[ 367] = 1'b1; frame1.error[ 367] = 1'b0;frame1.data[ 368] = 8'h63; frame1.valid[ 368] = 1'b1; frame1.error[ 368] = 1'b0;frame1.data[ 369] = 8'h64; frame1.valid[ 369] = 1'b1; frame1.error[ 369] = 1'b0;frame1.data[ 370] = 8'h65; frame1.valid[ 370] = 1'b1; frame1.error[ 370] = 1'b0;frame1.data[ 371] = 8'h66; frame1.valid[ 371] = 1'b1; frame1.error[ 371] = 1'b0;frame1.data[ 372] = 8'h67; frame1.valid[ 372] = 1'b1; frame1.error[ 372] = 1'b0;frame1.data[ 373] = 8'h68; frame1.valid[ 373] = 1'b1; frame1.error[ 373] = 1'b0;frame1.data[ 374] = 8'h69; frame1.valid[ 374] = 1'b1; frame1.error[ 374] = 1'b0;frame1.data[ 375] = 8'h6A; frame1.valid[ 375] = 1'b1; frame1.error[ 375] = 1'b0;frame1.data[ 376] = 8'h6B; frame1.valid[ 376] = 1'b1; frame1.error[ 376] = 1'b0;frame1.data[ 377] = 8'h6C; frame1.valid[ 377] = 1'b1; frame1.error[ 377] = 1'b0;frame1.data[ 378] = 8'h6D; frame1.valid[ 378] = 1'b1; frame1.error[ 378] = 1'b0;frame1.data[ 379] = 8'h6E; frame1.valid[ 379] = 1'b1; frame1.error[ 379] = 1'b0;frame1.data[ 380] = 8'h6F; frame1.valid[ 380] = 1'b1; frame1.error[ 380] = 1'b0;frame1.data[ 381] = 8'h70; frame1.valid[ 381] = 1'b1; frame1.error[ 381] = 1'b0;
        frame1.data[ 382] = 8'h71; frame1.valid[ 382] = 1'b1; frame1.error[ 382] = 1'b0;frame1.data[ 383] = 8'h72; frame1.valid[ 383] = 1'b1; frame1.error[ 383] = 1'b0;frame1.data[ 384] = 8'h73; frame1.valid[ 384] = 1'b1; frame1.error[ 384] = 1'b0;frame1.data[ 385] = 8'h74; frame1.valid[ 385] = 1'b1; frame1.error[ 385] = 1'b0;frame1.data[ 386] = 8'h75; frame1.valid[ 386] = 1'b1; frame1.error[ 386] = 1'b0;frame1.data[ 387] = 8'h76; frame1.valid[ 387] = 1'b1; frame1.error[ 387] = 1'b0;frame1.data[ 388] = 8'h77; frame1.valid[ 388] = 1'b1; frame1.error[ 388] = 1'b0;frame1.data[ 389] = 8'h78; frame1.valid[ 389] = 1'b1; frame1.error[ 389] = 1'b0;frame1.data[ 390] = 8'h79; frame1.valid[ 390] = 1'b1; frame1.error[ 390] = 1'b0;frame1.data[ 391] = 8'h7A; frame1.valid[ 391] = 1'b1; frame1.error[ 391] = 1'b0;frame1.data[ 392] = 8'h7B; frame1.valid[ 392] = 1'b1; frame1.error[ 392] = 1'b0;frame1.data[ 393] = 8'h7C; frame1.valid[ 393] = 1'b1; frame1.error[ 393] = 1'b0;frame1.data[ 394] = 8'h7D; frame1.valid[ 394] = 1'b1; frame1.error[ 394] = 1'b0;frame1.data[ 395] = 8'h7E; frame1.valid[ 395] = 1'b1; frame1.error[ 395] = 1'b0;frame1.data[ 396] = 8'h7F; frame1.valid[ 396] = 1'b1; frame1.error[ 396] = 1'b0;frame1.data[ 397] = 8'h80; frame1.valid[ 397] = 1'b1; frame1.error[ 397] = 1'b0;
        frame1.data[ 398] = 8'h81; frame1.valid[ 398] = 1'b1; frame1.error[ 398] = 1'b0;frame1.data[ 399] = 8'h82; frame1.valid[ 399] = 1'b1; frame1.error[ 399] = 1'b0;frame1.data[ 400] = 8'h83; frame1.valid[ 400] = 1'b1; frame1.error[ 400] = 1'b0;frame1.data[ 401] = 8'h84; frame1.valid[ 401] = 1'b1; frame1.error[ 401] = 1'b0;frame1.data[ 402] = 8'h85; frame1.valid[ 402] = 1'b1; frame1.error[ 402] = 1'b0;frame1.data[ 403] = 8'h86; frame1.valid[ 403] = 1'b1; frame1.error[ 403] = 1'b0;frame1.data[ 404] = 8'h87; frame1.valid[ 404] = 1'b1; frame1.error[ 404] = 1'b0;frame1.data[ 405] = 8'h88; frame1.valid[ 405] = 1'b1; frame1.error[ 405] = 1'b0;frame1.data[ 406] = 8'h89; frame1.valid[ 406] = 1'b1; frame1.error[ 406] = 1'b0;frame1.data[ 407] = 8'h8A; frame1.valid[ 407] = 1'b1; frame1.error[ 407] = 1'b0;frame1.data[ 408] = 8'h8B; frame1.valid[ 408] = 1'b1; frame1.error[ 408] = 1'b0;frame1.data[ 409] = 8'h8C; frame1.valid[ 409] = 1'b1; frame1.error[ 409] = 1'b0;frame1.data[ 410] = 8'h8D; frame1.valid[ 410] = 1'b1; frame1.error[ 410] = 1'b0;frame1.data[ 411] = 8'h8E; frame1.valid[ 411] = 1'b1; frame1.error[ 411] = 1'b0;frame1.data[ 412] = 8'h8F; frame1.valid[ 412] = 1'b1; frame1.error[ 412] = 1'b0;frame1.data[ 413] = 8'h90; frame1.valid[ 413] = 1'b1; frame1.error[ 413] = 1'b0;
        frame1.data[ 414] = 8'h91; frame1.valid[ 414] = 1'b1; frame1.error[ 414] = 1'b0;frame1.data[ 415] = 8'h92; frame1.valid[ 415] = 1'b1; frame1.error[ 415] = 1'b0;frame1.data[ 416] = 8'h93; frame1.valid[ 416] = 1'b1; frame1.error[ 416] = 1'b0;frame1.data[ 417] = 8'h94; frame1.valid[ 417] = 1'b1; frame1.error[ 417] = 1'b0;frame1.data[ 418] = 8'h95; frame1.valid[ 418] = 1'b1; frame1.error[ 418] = 1'b0;frame1.data[ 419] = 8'h96; frame1.valid[ 419] = 1'b1; frame1.error[ 419] = 1'b0;frame1.data[ 420] = 8'h97; frame1.valid[ 420] = 1'b1; frame1.error[ 420] = 1'b0;frame1.data[ 421] = 8'h98; frame1.valid[ 421] = 1'b1; frame1.error[ 421] = 1'b0;frame1.data[ 422] = 8'h99; frame1.valid[ 422] = 1'b1; frame1.error[ 422] = 1'b0;frame1.data[ 423] = 8'h9A; frame1.valid[ 423] = 1'b1; frame1.error[ 423] = 1'b0;frame1.data[ 424] = 8'h9B; frame1.valid[ 424] = 1'b1; frame1.error[ 424] = 1'b0;frame1.data[ 425] = 8'h9C; frame1.valid[ 425] = 1'b1; frame1.error[ 425] = 1'b0;frame1.data[ 426] = 8'h9D; frame1.valid[ 426] = 1'b1; frame1.error[ 426] = 1'b0;frame1.data[ 427] = 8'h9E; frame1.valid[ 427] = 1'b1; frame1.error[ 427] = 1'b0;frame1.data[ 428] = 8'h9F; frame1.valid[ 428] = 1'b1; frame1.error[ 428] = 1'b0;frame1.data[ 429] = 8'hA0; frame1.valid[ 429] = 1'b1; frame1.error[ 429] = 1'b0;
        frame1.data[ 430] = 8'hA1; frame1.valid[ 430] = 1'b1; frame1.error[ 430] = 1'b0;frame1.data[ 431] = 8'hA2; frame1.valid[ 431] = 1'b1; frame1.error[ 431] = 1'b0;frame1.data[ 432] = 8'hA3; frame1.valid[ 432] = 1'b1; frame1.error[ 432] = 1'b0;frame1.data[ 433] = 8'hA4; frame1.valid[ 433] = 1'b1; frame1.error[ 433] = 1'b0;frame1.data[ 434] = 8'hA5; frame1.valid[ 434] = 1'b1; frame1.error[ 434] = 1'b0;frame1.data[ 435] = 8'hA6; frame1.valid[ 435] = 1'b1; frame1.error[ 435] = 1'b0;frame1.data[ 436] = 8'hA7; frame1.valid[ 436] = 1'b1; frame1.error[ 436] = 1'b0;frame1.data[ 437] = 8'hA8; frame1.valid[ 437] = 1'b1; frame1.error[ 437] = 1'b0;frame1.data[ 438] = 8'hA9; frame1.valid[ 438] = 1'b1; frame1.error[ 438] = 1'b0;frame1.data[ 439] = 8'hAA; frame1.valid[ 439] = 1'b1; frame1.error[ 439] = 1'b0;frame1.data[ 440] = 8'hAB; frame1.valid[ 440] = 1'b1; frame1.error[ 440] = 1'b0;frame1.data[ 441] = 8'hAC; frame1.valid[ 441] = 1'b1; frame1.error[ 441] = 1'b0;frame1.data[ 442] = 8'hAD; frame1.valid[ 442] = 1'b1; frame1.error[ 442] = 1'b0;frame1.data[ 443] = 8'hAE; frame1.valid[ 443] = 1'b1; frame1.error[ 443] = 1'b0;frame1.data[ 444] = 8'hAF; frame1.valid[ 444] = 1'b1; frame1.error[ 444] = 1'b0;frame1.data[ 445] = 8'hB0; frame1.valid[ 445] = 1'b1; frame1.error[ 445] = 1'b0;
        frame1.data[ 446] = 8'hB1; frame1.valid[ 446] = 1'b1; frame1.error[ 446] = 1'b0;frame1.data[ 447] = 8'hB2; frame1.valid[ 447] = 1'b1; frame1.error[ 447] = 1'b0;frame1.data[ 448] = 8'hB3; frame1.valid[ 448] = 1'b1; frame1.error[ 448] = 1'b0;frame1.data[ 449] = 8'hB4; frame1.valid[ 449] = 1'b1; frame1.error[ 449] = 1'b0;frame1.data[ 450] = 8'hB5; frame1.valid[ 450] = 1'b1; frame1.error[ 450] = 1'b0;frame1.data[ 451] = 8'hB6; frame1.valid[ 451] = 1'b1; frame1.error[ 451] = 1'b0;frame1.data[ 452] = 8'hB7; frame1.valid[ 452] = 1'b1; frame1.error[ 452] = 1'b0;frame1.data[ 453] = 8'hB8; frame1.valid[ 453] = 1'b1; frame1.error[ 453] = 1'b0;frame1.data[ 454] = 8'hB9; frame1.valid[ 454] = 1'b1; frame1.error[ 454] = 1'b0;frame1.data[ 455] = 8'hBA; frame1.valid[ 455] = 1'b1; frame1.error[ 455] = 1'b0;frame1.data[ 456] = 8'hBB; frame1.valid[ 456] = 1'b1; frame1.error[ 456] = 1'b0;frame1.data[ 457] = 8'hBC; frame1.valid[ 457] = 1'b1; frame1.error[ 457] = 1'b0;frame1.data[ 458] = 8'hBD; frame1.valid[ 458] = 1'b1; frame1.error[ 458] = 1'b0;frame1.data[ 459] = 8'hBE; frame1.valid[ 459] = 1'b1; frame1.error[ 459] = 1'b0;frame1.data[ 460] = 8'hBF; frame1.valid[ 460] = 1'b1; frame1.error[ 460] = 1'b0;frame1.data[ 461] = 8'hC0; frame1.valid[ 461] = 1'b1; frame1.error[ 461] = 1'b0;
        frame1.data[ 462] = 8'hC1; frame1.valid[ 462] = 1'b1; frame1.error[ 462] = 1'b0;frame1.data[ 463] = 8'hC2; frame1.valid[ 463] = 1'b1; frame1.error[ 463] = 1'b0;frame1.data[ 464] = 8'hC3; frame1.valid[ 464] = 1'b1; frame1.error[ 464] = 1'b0;frame1.data[ 465] = 8'hC4; frame1.valid[ 465] = 1'b1; frame1.error[ 465] = 1'b0;frame1.data[ 466] = 8'hC5; frame1.valid[ 466] = 1'b1; frame1.error[ 466] = 1'b0;frame1.data[ 467] = 8'hC6; frame1.valid[ 467] = 1'b1; frame1.error[ 467] = 1'b0;frame1.data[ 468] = 8'hC7; frame1.valid[ 468] = 1'b1; frame1.error[ 468] = 1'b0;frame1.data[ 469] = 8'hC8; frame1.valid[ 469] = 1'b1; frame1.error[ 469] = 1'b0;frame1.data[ 470] = 8'hC9; frame1.valid[ 470] = 1'b1; frame1.error[ 470] = 1'b0;frame1.data[ 471] = 8'hCA; frame1.valid[ 471] = 1'b1; frame1.error[ 471] = 1'b0;frame1.data[ 472] = 8'hCB; frame1.valid[ 472] = 1'b1; frame1.error[ 472] = 1'b0;frame1.data[ 473] = 8'hCC; frame1.valid[ 473] = 1'b1; frame1.error[ 473] = 1'b0;frame1.data[ 474] = 8'hCD; frame1.valid[ 474] = 1'b1; frame1.error[ 474] = 1'b0;frame1.data[ 475] = 8'hCE; frame1.valid[ 475] = 1'b1; frame1.error[ 475] = 1'b0;frame1.data[ 476] = 8'hCF; frame1.valid[ 476] = 1'b1; frame1.error[ 476] = 1'b0;frame1.data[ 477] = 8'hD0; frame1.valid[ 477] = 1'b1; frame1.error[ 477] = 1'b0;
        frame1.data[ 478] = 8'hD1; frame1.valid[ 478] = 1'b1; frame1.error[ 478] = 1'b0;frame1.data[ 479] = 8'hD2; frame1.valid[ 479] = 1'b1; frame1.error[ 479] = 1'b0;frame1.data[ 480] = 8'hD3; frame1.valid[ 480] = 1'b1; frame1.error[ 480] = 1'b0;frame1.data[ 481] = 8'hD4; frame1.valid[ 481] = 1'b1; frame1.error[ 481] = 1'b0;frame1.data[ 482] = 8'hD5; frame1.valid[ 482] = 1'b1; frame1.error[ 482] = 1'b0;frame1.data[ 483] = 8'hD6; frame1.valid[ 483] = 1'b1; frame1.error[ 483] = 1'b0;frame1.data[ 484] = 8'hD7; frame1.valid[ 484] = 1'b1; frame1.error[ 484] = 1'b0;frame1.data[ 485] = 8'hD8; frame1.valid[ 485] = 1'b1; frame1.error[ 485] = 1'b0;frame1.data[ 486] = 8'hD9; frame1.valid[ 486] = 1'b1; frame1.error[ 486] = 1'b0;frame1.data[ 487] = 8'hDA; frame1.valid[ 487] = 1'b1; frame1.error[ 487] = 1'b0;frame1.data[ 488] = 8'hDB; frame1.valid[ 488] = 1'b1; frame1.error[ 488] = 1'b0;frame1.data[ 489] = 8'hDC; frame1.valid[ 489] = 1'b1; frame1.error[ 489] = 1'b0;frame1.data[ 490] = 8'hDD; frame1.valid[ 490] = 1'b1; frame1.error[ 490] = 1'b0;frame1.data[ 491] = 8'hDE; frame1.valid[ 491] = 1'b1; frame1.error[ 491] = 1'b0;frame1.data[ 492] = 8'hDF; frame1.valid[ 492] = 1'b1; frame1.error[ 492] = 1'b0;frame1.data[ 493] = 8'hE0; frame1.valid[ 493] = 1'b1; frame1.error[ 493] = 1'b0;
        frame1.data[ 494] = 8'hE1; frame1.valid[ 494] = 1'b1; frame1.error[ 494] = 1'b0;frame1.data[ 495] = 8'hE2; frame1.valid[ 495] = 1'b1; frame1.error[ 495] = 1'b0;frame1.data[ 496] = 8'hE3; frame1.valid[ 496] = 1'b1; frame1.error[ 496] = 1'b0;frame1.data[ 497] = 8'hE4; frame1.valid[ 497] = 1'b1; frame1.error[ 497] = 1'b0;frame1.data[ 498] = 8'hE5; frame1.valid[ 498] = 1'b1; frame1.error[ 498] = 1'b0;frame1.data[ 499] = 8'hE6; frame1.valid[ 499] = 1'b1; frame1.error[ 499] = 1'b0;frame1.data[ 500] = 8'hE7; frame1.valid[ 500] = 1'b1; frame1.error[ 500] = 1'b0;frame1.data[ 501] = 8'hE8; frame1.valid[ 501] = 1'b1; frame1.error[ 501] = 1'b0;frame1.data[ 502] = 8'hE9; frame1.valid[ 502] = 1'b1; frame1.error[ 502] = 1'b0;frame1.data[ 503] = 8'hEA; frame1.valid[ 503] = 1'b1; frame1.error[ 503] = 1'b0;frame1.data[ 504] = 8'hEB; frame1.valid[ 504] = 1'b1; frame1.error[ 504] = 1'b0;frame1.data[ 505] = 8'hEC; frame1.valid[ 505] = 1'b1; frame1.error[ 505] = 1'b0;frame1.data[ 506] = 8'hED; frame1.valid[ 506] = 1'b1; frame1.error[ 506] = 1'b0;frame1.data[ 507] = 8'hEE; frame1.valid[ 507] = 1'b1; frame1.error[ 507] = 1'b0;frame1.data[ 508] = 8'hEF; frame1.valid[ 508] = 1'b1; frame1.error[ 508] = 1'b0;frame1.data[ 509] = 8'hF0; frame1.valid[ 509] = 1'b1; frame1.error[ 509] = 1'b0;
        frame1.data[ 510] = 8'hF1; frame1.valid[ 510] = 1'b1; frame1.error[ 510] = 1'b0;frame1.data[ 511] = 8'hF2; frame1.valid[ 511] = 1'b1; frame1.error[ 511] = 1'b0;frame1.data[ 512] = 8'hF3; frame1.valid[ 512] = 1'b1; frame1.error[ 512] = 1'b0;frame1.data[ 513] = 8'hF4; frame1.valid[ 513] = 1'b1; frame1.error[ 513] = 1'b0;frame1.data[ 514] = 8'hF5; frame1.valid[ 514] = 1'b1; frame1.error[ 514] = 1'b0;frame1.data[ 515] = 8'hF6; frame1.valid[ 515] = 1'b1; frame1.error[ 515] = 1'b0;frame1.data[ 516] = 8'hF7; frame1.valid[ 516] = 1'b1; frame1.error[ 516] = 1'b0;frame1.data[ 517] = 8'hF8; frame1.valid[ 517] = 1'b1; frame1.error[ 517] = 1'b0;frame1.data[ 518] = 8'hF9; frame1.valid[ 518] = 1'b1; frame1.error[ 518] = 1'b0;frame1.data[ 519] = 8'hFA; frame1.valid[ 519] = 1'b1; frame1.error[ 519] = 1'b0;frame1.data[ 520] = 8'hFB; frame1.valid[ 520] = 1'b1; frame1.error[ 520] = 1'b0;frame1.data[ 521] = 8'hFC; frame1.valid[ 521] = 1'b1; frame1.error[ 521] = 1'b0;frame1.data[ 522] = 8'hFD; frame1.valid[ 522] = 1'b1; frame1.error[ 522] = 1'b0;frame1.data[ 523] = 8'hFE; frame1.valid[ 523] = 1'b1; frame1.error[ 523] = 1'b0;frame1.data[ 524] = 8'h00; frame1.valid[ 524] = 1'b1; frame1.error[ 524] = 1'b0;frame1.data[ 525] = 8'h01; frame1.valid[ 525] = 1'b1; frame1.error[ 525] = 1'b0;
        frame1.data[ 526] = 8'h02; frame1.valid[ 526] = 1'b1; frame1.error[ 526] = 1'b0;frame1.data[ 527] = 8'h03; frame1.valid[ 527] = 1'b1; frame1.error[ 527] = 1'b0;frame1.data[ 528] = 8'h04; frame1.valid[ 528] = 1'b1; frame1.error[ 528] = 1'b0;frame1.data[ 529] = 8'h05; frame1.valid[ 529] = 1'b1; frame1.error[ 529] = 1'b0;frame1.data[ 530] = 8'h06; frame1.valid[ 530] = 1'b1; frame1.error[ 530] = 1'b0;frame1.data[ 531] = 8'h07; frame1.valid[ 531] = 1'b1; frame1.error[ 531] = 1'b0;frame1.data[ 532] = 8'h08; frame1.valid[ 532] = 1'b1; frame1.error[ 532] = 1'b0;frame1.data[ 533] = 8'h09; frame1.valid[ 533] = 1'b1; frame1.error[ 533] = 1'b0;frame1.data[ 534] = 8'h0A; frame1.valid[ 534] = 1'b1; frame1.error[ 534] = 1'b0;frame1.data[ 535] = 8'h0B; frame1.valid[ 535] = 1'b1; frame1.error[ 535] = 1'b0;frame1.data[ 536] = 8'h0C; frame1.valid[ 536] = 1'b1; frame1.error[ 536] = 1'b0;frame1.data[ 537] = 8'h0D; frame1.valid[ 537] = 1'b1; frame1.error[ 537] = 1'b0;frame1.data[ 538] = 8'h0E; frame1.valid[ 538] = 1'b1; frame1.error[ 538] = 1'b0;frame1.data[ 539] = 8'h0F; frame1.valid[ 539] = 1'b1; frame1.error[ 539] = 1'b0;frame1.data[ 540] = 8'h10; frame1.valid[ 540] = 1'b1; frame1.error[ 540] = 1'b0;frame1.data[ 541] = 8'h11; frame1.valid[ 541] = 1'b1; frame1.error[ 541] = 1'b0;
        frame1.data[ 542] = 8'h12; frame1.valid[ 542] = 1'b1; frame1.error[ 542] = 1'b0;frame1.data[ 543] = 8'h13; frame1.valid[ 543] = 1'b1; frame1.error[ 543] = 1'b0;frame1.data[ 544] = 8'h14; frame1.valid[ 544] = 1'b1; frame1.error[ 544] = 1'b0;frame1.data[ 545] = 8'h15; frame1.valid[ 545] = 1'b1; frame1.error[ 545] = 1'b0;frame1.data[ 546] = 8'h16; frame1.valid[ 546] = 1'b1; frame1.error[ 546] = 1'b0;frame1.data[ 547] = 8'h17; frame1.valid[ 547] = 1'b1; frame1.error[ 547] = 1'b0;frame1.data[ 548] = 8'h18; frame1.valid[ 548] = 1'b1; frame1.error[ 548] = 1'b0;frame1.data[ 549] = 8'h19; frame1.valid[ 549] = 1'b1; frame1.error[ 549] = 1'b0;frame1.data[ 550] = 8'h1A; frame1.valid[ 550] = 1'b1; frame1.error[ 550] = 1'b0;frame1.data[ 551] = 8'h1B; frame1.valid[ 551] = 1'b1; frame1.error[ 551] = 1'b0;frame1.data[ 552] = 8'h1C; frame1.valid[ 552] = 1'b1; frame1.error[ 552] = 1'b0;frame1.data[ 553] = 8'h1D; frame1.valid[ 553] = 1'b1; frame1.error[ 553] = 1'b0;frame1.data[ 554] = 8'h1E; frame1.valid[ 554] = 1'b1; frame1.error[ 554] = 1'b0;frame1.data[ 555] = 8'h1F; frame1.valid[ 555] = 1'b1; frame1.error[ 555] = 1'b0;frame1.data[ 556] = 8'h20; frame1.valid[ 556] = 1'b1; frame1.error[ 556] = 1'b0;frame1.data[ 557] = 8'h21; frame1.valid[ 557] = 1'b1; frame1.error[ 557] = 1'b0;
        frame1.data[ 558] = 8'h22; frame1.valid[ 558] = 1'b1; frame1.error[ 558] = 1'b0;frame1.data[ 559] = 8'h23; frame1.valid[ 559] = 1'b1; frame1.error[ 559] = 1'b0;frame1.data[ 560] = 8'h24; frame1.valid[ 560] = 1'b1; frame1.error[ 560] = 1'b0;frame1.data[ 561] = 8'h25; frame1.valid[ 561] = 1'b1; frame1.error[ 561] = 1'b0;frame1.data[ 562] = 8'h26; frame1.valid[ 562] = 1'b1; frame1.error[ 562] = 1'b0;frame1.data[ 563] = 8'h27; frame1.valid[ 563] = 1'b1; frame1.error[ 563] = 1'b0;frame1.data[ 564] = 8'h28; frame1.valid[ 564] = 1'b1; frame1.error[ 564] = 1'b0;frame1.data[ 565] = 8'h29; frame1.valid[ 565] = 1'b1; frame1.error[ 565] = 1'b0;frame1.data[ 566] = 8'h2A; frame1.valid[ 566] = 1'b1; frame1.error[ 566] = 1'b0;frame1.data[ 567] = 8'h2B; frame1.valid[ 567] = 1'b1; frame1.error[ 567] = 1'b0;frame1.data[ 568] = 8'h2C; frame1.valid[ 568] = 1'b1; frame1.error[ 568] = 1'b0;frame1.data[ 569] = 8'h2D; frame1.valid[ 569] = 1'b1; frame1.error[ 569] = 1'b0;frame1.data[ 570] = 8'h2E; frame1.valid[ 570] = 1'b1; frame1.error[ 570] = 1'b0;frame1.data[ 571] = 8'h2F; frame1.valid[ 571] = 1'b1; frame1.error[ 571] = 1'b0;frame1.data[ 572] = 8'h30; frame1.valid[ 572] = 1'b1; frame1.error[ 572] = 1'b0;frame1.data[ 573] = 8'h31; frame1.valid[ 573] = 1'b1; frame1.error[ 573] = 1'b0;
        frame1.data[ 574] = 8'h32; frame1.valid[ 574] = 1'b1; frame1.error[ 574] = 1'b0;frame1.data[ 575] = 8'h33; frame1.valid[ 575] = 1'b1; frame1.error[ 575] = 1'b0;frame1.data[ 576] = 8'h34; frame1.valid[ 576] = 1'b1; frame1.error[ 576] = 1'b0;frame1.data[ 577] = 8'h35; frame1.valid[ 577] = 1'b1; frame1.error[ 577] = 1'b0;frame1.data[ 578] = 8'h36; frame1.valid[ 578] = 1'b1; frame1.error[ 578] = 1'b0;frame1.data[ 579] = 8'h37; frame1.valid[ 579] = 1'b1; frame1.error[ 579] = 1'b0;frame1.data[ 580] = 8'h38; frame1.valid[ 580] = 1'b1; frame1.error[ 580] = 1'b0;frame1.data[ 581] = 8'h39; frame1.valid[ 581] = 1'b1; frame1.error[ 581] = 1'b0;frame1.data[ 582] = 8'h3A; frame1.valid[ 582] = 1'b1; frame1.error[ 582] = 1'b0;frame1.data[ 583] = 8'h3B; frame1.valid[ 583] = 1'b1; frame1.error[ 583] = 1'b0;frame1.data[ 584] = 8'h3C; frame1.valid[ 584] = 1'b1; frame1.error[ 584] = 1'b0;frame1.data[ 585] = 8'h3D; frame1.valid[ 585] = 1'b1; frame1.error[ 585] = 1'b0;frame1.data[ 586] = 8'h3E; frame1.valid[ 586] = 1'b1; frame1.error[ 586] = 1'b0;frame1.data[ 587] = 8'h3F; frame1.valid[ 587] = 1'b1; frame1.error[ 587] = 1'b0;frame1.data[ 588] = 8'h40; frame1.valid[ 588] = 1'b1; frame1.error[ 588] = 1'b0;frame1.data[ 589] = 8'h41; frame1.valid[ 589] = 1'b1; frame1.error[ 589] = 1'b0;
        frame1.data[ 590] = 8'h42; frame1.valid[ 590] = 1'b1; frame1.error[ 590] = 1'b0;frame1.data[ 591] = 8'h43; frame1.valid[ 591] = 1'b1; frame1.error[ 591] = 1'b0;frame1.data[ 592] = 8'h44; frame1.valid[ 592] = 1'b1; frame1.error[ 592] = 1'b0;frame1.data[ 593] = 8'h45; frame1.valid[ 593] = 1'b1; frame1.error[ 593] = 1'b0;frame1.data[ 594] = 8'h46; frame1.valid[ 594] = 1'b1; frame1.error[ 594] = 1'b0;frame1.data[ 595] = 8'h47; frame1.valid[ 595] = 1'b1; frame1.error[ 595] = 1'b0;frame1.data[ 596] = 8'h48; frame1.valid[ 596] = 1'b1; frame1.error[ 596] = 1'b0;frame1.data[ 597] = 8'h49; frame1.valid[ 597] = 1'b1; frame1.error[ 597] = 1'b0;frame1.data[ 598] = 8'h4A; frame1.valid[ 598] = 1'b1; frame1.error[ 598] = 1'b0;frame1.data[ 599] = 8'h4B; frame1.valid[ 599] = 1'b1; frame1.error[ 599] = 1'b0;frame1.data[ 600] = 8'h4C; frame1.valid[ 600] = 1'b1; frame1.error[ 600] = 1'b0;frame1.data[ 601] = 8'h4D; frame1.valid[ 601] = 1'b1; frame1.error[ 601] = 1'b0;frame1.data[ 602] = 8'h4E; frame1.valid[ 602] = 1'b1; frame1.error[ 602] = 1'b0;frame1.data[ 603] = 8'h4F; frame1.valid[ 603] = 1'b1; frame1.error[ 603] = 1'b0;frame1.data[ 604] = 8'h50; frame1.valid[ 604] = 1'b1; frame1.error[ 604] = 1'b0;frame1.data[ 605] = 8'h51; frame1.valid[ 605] = 1'b1; frame1.error[ 605] = 1'b0;
        frame1.data[ 606] = 8'h52; frame1.valid[ 606] = 1'b1; frame1.error[ 606] = 1'b0;frame1.data[ 607] = 8'h53; frame1.valid[ 607] = 1'b1; frame1.error[ 607] = 1'b0;frame1.data[ 608] = 8'h54; frame1.valid[ 608] = 1'b1; frame1.error[ 608] = 1'b0;frame1.data[ 609] = 8'h55; frame1.valid[ 609] = 1'b1; frame1.error[ 609] = 1'b0;frame1.data[ 610] = 8'h56; frame1.valid[ 610] = 1'b1; frame1.error[ 610] = 1'b0;frame1.data[ 611] = 8'h57; frame1.valid[ 611] = 1'b1; frame1.error[ 611] = 1'b0;frame1.data[ 612] = 8'h58; frame1.valid[ 612] = 1'b1; frame1.error[ 612] = 1'b0;frame1.data[ 613] = 8'h59; frame1.valid[ 613] = 1'b1; frame1.error[ 613] = 1'b0;frame1.data[ 614] = 8'h5A; frame1.valid[ 614] = 1'b1; frame1.error[ 614] = 1'b0;frame1.data[ 615] = 8'h5B; frame1.valid[ 615] = 1'b1; frame1.error[ 615] = 1'b0;frame1.data[ 616] = 8'h5C; frame1.valid[ 616] = 1'b1; frame1.error[ 616] = 1'b0;frame1.data[ 617] = 8'h5D; frame1.valid[ 617] = 1'b1; frame1.error[ 617] = 1'b0;frame1.data[ 618] = 8'h5E; frame1.valid[ 618] = 1'b1; frame1.error[ 618] = 1'b0;frame1.data[ 619] = 8'h5F; frame1.valid[ 619] = 1'b1; frame1.error[ 619] = 1'b0;frame1.data[ 620] = 8'h60; frame1.valid[ 620] = 1'b1; frame1.error[ 620] = 1'b0;frame1.data[ 621] = 8'h61; frame1.valid[ 621] = 1'b1; frame1.error[ 621] = 1'b0;
        frame1.data[ 622] = 8'h62; frame1.valid[ 622] = 1'b1; frame1.error[ 622] = 1'b0;frame1.data[ 623] = 8'h63; frame1.valid[ 623] = 1'b1; frame1.error[ 623] = 1'b0;frame1.data[ 624] = 8'h64; frame1.valid[ 624] = 1'b1; frame1.error[ 624] = 1'b0;frame1.data[ 625] = 8'h65; frame1.valid[ 625] = 1'b1; frame1.error[ 625] = 1'b0;frame1.data[ 626] = 8'h66; frame1.valid[ 626] = 1'b1; frame1.error[ 626] = 1'b0;frame1.data[ 627] = 8'h67; frame1.valid[ 627] = 1'b1; frame1.error[ 627] = 1'b0;frame1.data[ 628] = 8'h68; frame1.valid[ 628] = 1'b1; frame1.error[ 628] = 1'b0;frame1.data[ 629] = 8'h69; frame1.valid[ 629] = 1'b1; frame1.error[ 629] = 1'b0;frame1.data[ 630] = 8'h6A; frame1.valid[ 630] = 1'b1; frame1.error[ 630] = 1'b0;frame1.data[ 631] = 8'h6B; frame1.valid[ 631] = 1'b1; frame1.error[ 631] = 1'b0;frame1.data[ 632] = 8'h6C; frame1.valid[ 632] = 1'b1; frame1.error[ 632] = 1'b0;frame1.data[ 633] = 8'h6D; frame1.valid[ 633] = 1'b1; frame1.error[ 633] = 1'b0;frame1.data[ 634] = 8'h6E; frame1.valid[ 634] = 1'b1; frame1.error[ 634] = 1'b0;frame1.data[ 635] = 8'h6F; frame1.valid[ 635] = 1'b1; frame1.error[ 635] = 1'b0;frame1.data[ 636] = 8'h70; frame1.valid[ 636] = 1'b1; frame1.error[ 636] = 1'b0;frame1.data[ 637] = 8'h71; frame1.valid[ 637] = 1'b1; frame1.error[ 637] = 1'b0;
        frame1.data[ 638] = 8'h72; frame1.valid[ 638] = 1'b1; frame1.error[ 638] = 1'b0;frame1.data[ 639] = 8'h73; frame1.valid[ 639] = 1'b1; frame1.error[ 639] = 1'b0;frame1.data[ 640] = 8'h74; frame1.valid[ 640] = 1'b1; frame1.error[ 640] = 1'b0;frame1.data[ 641] = 8'h75; frame1.valid[ 641] = 1'b1; frame1.error[ 641] = 1'b0;frame1.data[ 642] = 8'h76; frame1.valid[ 642] = 1'b1; frame1.error[ 642] = 1'b0;frame1.data[ 643] = 8'h77; frame1.valid[ 643] = 1'b1; frame1.error[ 643] = 1'b0;frame1.data[ 644] = 8'h78; frame1.valid[ 644] = 1'b1; frame1.error[ 644] = 1'b0;frame1.data[ 645] = 8'h79; frame1.valid[ 645] = 1'b1; frame1.error[ 645] = 1'b0;frame1.data[ 646] = 8'h7A; frame1.valid[ 646] = 1'b1; frame1.error[ 646] = 1'b0;frame1.data[ 647] = 8'h7B; frame1.valid[ 647] = 1'b1; frame1.error[ 647] = 1'b0;frame1.data[ 648] = 8'h7C; frame1.valid[ 648] = 1'b1; frame1.error[ 648] = 1'b0;frame1.data[ 649] = 8'h7D; frame1.valid[ 649] = 1'b1; frame1.error[ 649] = 1'b0;frame1.data[ 650] = 8'h7E; frame1.valid[ 650] = 1'b1; frame1.error[ 650] = 1'b0;frame1.data[ 651] = 8'h7F; frame1.valid[ 651] = 1'b1; frame1.error[ 651] = 1'b0;frame1.data[ 652] = 8'h80; frame1.valid[ 652] = 1'b1; frame1.error[ 652] = 1'b0;frame1.data[ 653] = 8'h81; frame1.valid[ 653] = 1'b1; frame1.error[ 653] = 1'b0;
        frame1.data[ 654] = 8'h82; frame1.valid[ 654] = 1'b1; frame1.error[ 654] = 1'b0;frame1.data[ 655] = 8'h83; frame1.valid[ 655] = 1'b1; frame1.error[ 655] = 1'b0;frame1.data[ 656] = 8'h84; frame1.valid[ 656] = 1'b1; frame1.error[ 656] = 1'b0;frame1.data[ 657] = 8'h85; frame1.valid[ 657] = 1'b1; frame1.error[ 657] = 1'b0;frame1.data[ 658] = 8'h86; frame1.valid[ 658] = 1'b1; frame1.error[ 658] = 1'b0;frame1.data[ 659] = 8'h87; frame1.valid[ 659] = 1'b1; frame1.error[ 659] = 1'b0;frame1.data[ 660] = 8'h88; frame1.valid[ 660] = 1'b1; frame1.error[ 660] = 1'b0;frame1.data[ 661] = 8'h89; frame1.valid[ 661] = 1'b1; frame1.error[ 661] = 1'b0;frame1.data[ 662] = 8'h8A; frame1.valid[ 662] = 1'b1; frame1.error[ 662] = 1'b0;frame1.data[ 663] = 8'h8B; frame1.valid[ 663] = 1'b1; frame1.error[ 663] = 1'b0;frame1.data[ 664] = 8'h8C; frame1.valid[ 664] = 1'b1; frame1.error[ 664] = 1'b0;frame1.data[ 665] = 8'h8D; frame1.valid[ 665] = 1'b1; frame1.error[ 665] = 1'b0;frame1.data[ 666] = 8'h8E; frame1.valid[ 666] = 1'b1; frame1.error[ 666] = 1'b0;frame1.data[ 667] = 8'h8F; frame1.valid[ 667] = 1'b1; frame1.error[ 667] = 1'b0;frame1.data[ 668] = 8'h90; frame1.valid[ 668] = 1'b1; frame1.error[ 668] = 1'b0;frame1.data[ 669] = 8'h91; frame1.valid[ 669] = 1'b1; frame1.error[ 669] = 1'b0;
        frame1.data[ 670] = 8'h92; frame1.valid[ 670] = 1'b1; frame1.error[ 670] = 1'b0;frame1.data[ 671] = 8'h93; frame1.valid[ 671] = 1'b1; frame1.error[ 671] = 1'b0;frame1.data[ 672] = 8'h94; frame1.valid[ 672] = 1'b1; frame1.error[ 672] = 1'b0;frame1.data[ 673] = 8'h95; frame1.valid[ 673] = 1'b1; frame1.error[ 673] = 1'b0;frame1.data[ 674] = 8'h96; frame1.valid[ 674] = 1'b1; frame1.error[ 674] = 1'b0;frame1.data[ 675] = 8'h97; frame1.valid[ 675] = 1'b1; frame1.error[ 675] = 1'b0;frame1.data[ 676] = 8'h98; frame1.valid[ 676] = 1'b1; frame1.error[ 676] = 1'b0;frame1.data[ 677] = 8'h99; frame1.valid[ 677] = 1'b1; frame1.error[ 677] = 1'b0;frame1.data[ 678] = 8'h9A; frame1.valid[ 678] = 1'b1; frame1.error[ 678] = 1'b0;frame1.data[ 679] = 8'h9B; frame1.valid[ 679] = 1'b1; frame1.error[ 679] = 1'b0;frame1.data[ 680] = 8'h9C; frame1.valid[ 680] = 1'b1; frame1.error[ 680] = 1'b0;frame1.data[ 681] = 8'h9D; frame1.valid[ 681] = 1'b1; frame1.error[ 681] = 1'b0;frame1.data[ 682] = 8'h9E; frame1.valid[ 682] = 1'b1; frame1.error[ 682] = 1'b0;frame1.data[ 683] = 8'h9F; frame1.valid[ 683] = 1'b1; frame1.error[ 683] = 1'b0;frame1.data[ 684] = 8'hA0; frame1.valid[ 684] = 1'b1; frame1.error[ 684] = 1'b0;frame1.data[ 685] = 8'hA1; frame1.valid[ 685] = 1'b1; frame1.error[ 685] = 1'b0;
        frame1.data[ 686] = 8'hA2; frame1.valid[ 686] = 1'b1; frame1.error[ 686] = 1'b0;frame1.data[ 687] = 8'hA3; frame1.valid[ 687] = 1'b1; frame1.error[ 687] = 1'b0;frame1.data[ 688] = 8'hA4; frame1.valid[ 688] = 1'b1; frame1.error[ 688] = 1'b0;frame1.data[ 689] = 8'hA5; frame1.valid[ 689] = 1'b1; frame1.error[ 689] = 1'b0;frame1.data[ 690] = 8'hA6; frame1.valid[ 690] = 1'b1; frame1.error[ 690] = 1'b0;frame1.data[ 691] = 8'hA7; frame1.valid[ 691] = 1'b1; frame1.error[ 691] = 1'b0;frame1.data[ 692] = 8'hA8; frame1.valid[ 692] = 1'b1; frame1.error[ 692] = 1'b0;frame1.data[ 693] = 8'hA9; frame1.valid[ 693] = 1'b1; frame1.error[ 693] = 1'b0;frame1.data[ 694] = 8'hAA; frame1.valid[ 694] = 1'b1; frame1.error[ 694] = 1'b0;frame1.data[ 695] = 8'hAB; frame1.valid[ 695] = 1'b1; frame1.error[ 695] = 1'b0;frame1.data[ 696] = 8'hAC; frame1.valid[ 696] = 1'b1; frame1.error[ 696] = 1'b0;frame1.data[ 697] = 8'hAD; frame1.valid[ 697] = 1'b1; frame1.error[ 697] = 1'b0;frame1.data[ 698] = 8'hAE; frame1.valid[ 698] = 1'b1; frame1.error[ 698] = 1'b0;frame1.data[ 699] = 8'hAF; frame1.valid[ 699] = 1'b1; frame1.error[ 699] = 1'b0;frame1.data[ 700] = 8'hB0; frame1.valid[ 700] = 1'b1; frame1.error[ 700] = 1'b0;frame1.data[ 701] = 8'hB1; frame1.valid[ 701] = 1'b1; frame1.error[ 701] = 1'b0;
        frame1.data[ 702] = 8'hB2; frame1.valid[ 702] = 1'b1; frame1.error[ 702] = 1'b0;frame1.data[ 703] = 8'hB3; frame1.valid[ 703] = 1'b1; frame1.error[ 703] = 1'b0;frame1.data[ 704] = 8'hB4; frame1.valid[ 704] = 1'b1; frame1.error[ 704] = 1'b0;frame1.data[ 705] = 8'hB5; frame1.valid[ 705] = 1'b1; frame1.error[ 705] = 1'b0;frame1.data[ 706] = 8'hB6; frame1.valid[ 706] = 1'b1; frame1.error[ 706] = 1'b0;frame1.data[ 707] = 8'hB7; frame1.valid[ 707] = 1'b1; frame1.error[ 707] = 1'b0;frame1.data[ 708] = 8'hB8; frame1.valid[ 708] = 1'b1; frame1.error[ 708] = 1'b0;frame1.data[ 709] = 8'hB9; frame1.valid[ 709] = 1'b1; frame1.error[ 709] = 1'b0;frame1.data[ 710] = 8'hBA; frame1.valid[ 710] = 1'b1; frame1.error[ 710] = 1'b0;frame1.data[ 711] = 8'hBB; frame1.valid[ 711] = 1'b1; frame1.error[ 711] = 1'b0;frame1.data[ 712] = 8'hBC; frame1.valid[ 712] = 1'b1; frame1.error[ 712] = 1'b0;frame1.data[ 713] = 8'hBD; frame1.valid[ 713] = 1'b1; frame1.error[ 713] = 1'b0;frame1.data[ 714] = 8'hBE; frame1.valid[ 714] = 1'b1; frame1.error[ 714] = 1'b0;frame1.data[ 715] = 8'hBF; frame1.valid[ 715] = 1'b1; frame1.error[ 715] = 1'b0;frame1.data[ 716] = 8'hC0; frame1.valid[ 716] = 1'b1; frame1.error[ 716] = 1'b0;frame1.data[ 717] = 8'hC1; frame1.valid[ 717] = 1'b1; frame1.error[ 717] = 1'b0;
        frame1.data[ 718] = 8'hC2; frame1.valid[ 718] = 1'b1; frame1.error[ 718] = 1'b0;frame1.data[ 719] = 8'hC3; frame1.valid[ 719] = 1'b1; frame1.error[ 719] = 1'b0;frame1.data[ 720] = 8'hC4; frame1.valid[ 720] = 1'b1; frame1.error[ 720] = 1'b0;frame1.data[ 721] = 8'hC5; frame1.valid[ 721] = 1'b1; frame1.error[ 721] = 1'b0;frame1.data[ 722] = 8'hC6; frame1.valid[ 722] = 1'b1; frame1.error[ 722] = 1'b0;frame1.data[ 723] = 8'hC7; frame1.valid[ 723] = 1'b1; frame1.error[ 723] = 1'b0;frame1.data[ 724] = 8'hC8; frame1.valid[ 724] = 1'b1; frame1.error[ 724] = 1'b0;frame1.data[ 725] = 8'hC9; frame1.valid[ 725] = 1'b1; frame1.error[ 725] = 1'b0;frame1.data[ 726] = 8'hCA; frame1.valid[ 726] = 1'b1; frame1.error[ 726] = 1'b0;frame1.data[ 727] = 8'hCB; frame1.valid[ 727] = 1'b1; frame1.error[ 727] = 1'b0;frame1.data[ 728] = 8'hCC; frame1.valid[ 728] = 1'b1; frame1.error[ 728] = 1'b0;frame1.data[ 729] = 8'hCD; frame1.valid[ 729] = 1'b1; frame1.error[ 729] = 1'b0;frame1.data[ 730] = 8'hCE; frame1.valid[ 730] = 1'b1; frame1.error[ 730] = 1'b0;frame1.data[ 731] = 8'hCF; frame1.valid[ 731] = 1'b1; frame1.error[ 731] = 1'b0;frame1.data[ 732] = 8'hD0; frame1.valid[ 732] = 1'b1; frame1.error[ 732] = 1'b0;frame1.data[ 733] = 8'hD1; frame1.valid[ 733] = 1'b1; frame1.error[ 733] = 1'b0;
        frame1.data[ 734] = 8'hD2; frame1.valid[ 734] = 1'b1; frame1.error[ 734] = 1'b0;frame1.data[ 735] = 8'hD3; frame1.valid[ 735] = 1'b1; frame1.error[ 735] = 1'b0;frame1.data[ 736] = 8'hD4; frame1.valid[ 736] = 1'b1; frame1.error[ 736] = 1'b0;frame1.data[ 737] = 8'hD5; frame1.valid[ 737] = 1'b1; frame1.error[ 737] = 1'b0;frame1.data[ 738] = 8'hD6; frame1.valid[ 738] = 1'b1; frame1.error[ 738] = 1'b0;frame1.data[ 739] = 8'hD7; frame1.valid[ 739] = 1'b1; frame1.error[ 739] = 1'b0;frame1.data[ 740] = 8'hD8; frame1.valid[ 740] = 1'b1; frame1.error[ 740] = 1'b0;frame1.data[ 741] = 8'hD9; frame1.valid[ 741] = 1'b1; frame1.error[ 741] = 1'b0;frame1.data[ 742] = 8'hDA; frame1.valid[ 742] = 1'b1; frame1.error[ 742] = 1'b0;frame1.data[ 743] = 8'hDB; frame1.valid[ 743] = 1'b1; frame1.error[ 743] = 1'b0;frame1.data[ 744] = 8'hDC; frame1.valid[ 744] = 1'b1; frame1.error[ 744] = 1'b0;frame1.data[ 745] = 8'hDD; frame1.valid[ 745] = 1'b1; frame1.error[ 745] = 1'b0;frame1.data[ 746] = 8'hDE; frame1.valid[ 746] = 1'b1; frame1.error[ 746] = 1'b0;frame1.data[ 747] = 8'hDF; frame1.valid[ 747] = 1'b1; frame1.error[ 747] = 1'b0;frame1.data[ 748] = 8'hE0; frame1.valid[ 748] = 1'b1; frame1.error[ 748] = 1'b0;frame1.data[ 749] = 8'hE1; frame1.valid[ 749] = 1'b1; frame1.error[ 749] = 1'b0;
        frame1.data[ 750] = 8'hE2; frame1.valid[ 750] = 1'b1; frame1.error[ 750] = 1'b0;frame1.data[ 751] = 8'hE3; frame1.valid[ 751] = 1'b1; frame1.error[ 751] = 1'b0;frame1.data[ 752] = 8'hE4; frame1.valid[ 752] = 1'b1; frame1.error[ 752] = 1'b0;frame1.data[ 753] = 8'hE5; frame1.valid[ 753] = 1'b1; frame1.error[ 753] = 1'b0;frame1.data[ 754] = 8'hE6; frame1.valid[ 754] = 1'b1; frame1.error[ 754] = 1'b0;frame1.data[ 755] = 8'hE7; frame1.valid[ 755] = 1'b1; frame1.error[ 755] = 1'b0;frame1.data[ 756] = 8'hE8; frame1.valid[ 756] = 1'b1; frame1.error[ 756] = 1'b0;frame1.data[ 757] = 8'hE9; frame1.valid[ 757] = 1'b1; frame1.error[ 757] = 1'b0;frame1.data[ 758] = 8'hEA; frame1.valid[ 758] = 1'b1; frame1.error[ 758] = 1'b0;frame1.data[ 759] = 8'hEB; frame1.valid[ 759] = 1'b1; frame1.error[ 759] = 1'b0;frame1.data[ 760] = 8'hEC; frame1.valid[ 760] = 1'b1; frame1.error[ 760] = 1'b0;frame1.data[ 761] = 8'hED; frame1.valid[ 761] = 1'b1; frame1.error[ 761] = 1'b0;frame1.data[ 762] = 8'hEE; frame1.valid[ 762] = 1'b1; frame1.error[ 762] = 1'b0;frame1.data[ 763] = 8'hEF; frame1.valid[ 763] = 1'b1; frame1.error[ 763] = 1'b0;frame1.data[ 764] = 8'hF0; frame1.valid[ 764] = 1'b1; frame1.error[ 764] = 1'b0;frame1.data[ 765] = 8'hF1; frame1.valid[ 765] = 1'b1; frame1.error[ 765] = 1'b0;
        frame1.data[ 766] = 8'hF2; frame1.valid[ 766] = 1'b1; frame1.error[ 766] = 1'b0;frame1.data[ 767] = 8'hF3; frame1.valid[ 767] = 1'b1; frame1.error[ 767] = 1'b0;frame1.data[ 768] = 8'hF4; frame1.valid[ 768] = 1'b1; frame1.error[ 768] = 1'b0;frame1.data[ 769] = 8'hF5; frame1.valid[ 769] = 1'b1; frame1.error[ 769] = 1'b0;frame1.data[ 770] = 8'hF6; frame1.valid[ 770] = 1'b1; frame1.error[ 770] = 1'b0;frame1.data[ 771] = 8'hF7; frame1.valid[ 771] = 1'b1; frame1.error[ 771] = 1'b0;frame1.data[ 772] = 8'hF8; frame1.valid[ 772] = 1'b1; frame1.error[ 772] = 1'b0;frame1.data[ 773] = 8'hF9; frame1.valid[ 773] = 1'b1; frame1.error[ 773] = 1'b0;frame1.data[ 774] = 8'hFA; frame1.valid[ 774] = 1'b1; frame1.error[ 774] = 1'b0;frame1.data[ 775] = 8'hFB; frame1.valid[ 775] = 1'b1; frame1.error[ 775] = 1'b0;frame1.data[ 776] = 8'hFC; frame1.valid[ 776] = 1'b1; frame1.error[ 776] = 1'b0;frame1.data[ 777] = 8'hFD; frame1.valid[ 777] = 1'b1; frame1.error[ 777] = 1'b0;frame1.data[ 778] = 8'hFE; frame1.valid[ 778] = 1'b1; frame1.error[ 778] = 1'b0;frame1.data[ 779] = 8'h00; frame1.valid[ 779] = 1'b1; frame1.error[ 779] = 1'b0;frame1.data[ 780] = 8'h01; frame1.valid[ 780] = 1'b1; frame1.error[ 780] = 1'b0;frame1.data[ 781] = 8'h02; frame1.valid[ 781] = 1'b1; frame1.error[ 781] = 1'b0;
        frame1.data[ 782] = 8'h03; frame1.valid[ 782] = 1'b1; frame1.error[ 782] = 1'b0;frame1.data[ 783] = 8'h04; frame1.valid[ 783] = 1'b1; frame1.error[ 783] = 1'b0;frame1.data[ 784] = 8'h05; frame1.valid[ 784] = 1'b1; frame1.error[ 784] = 1'b0;frame1.data[ 785] = 8'h06; frame1.valid[ 785] = 1'b1; frame1.error[ 785] = 1'b0;frame1.data[ 786] = 8'h07; frame1.valid[ 786] = 1'b1; frame1.error[ 786] = 1'b0;frame1.data[ 787] = 8'h08; frame1.valid[ 787] = 1'b1; frame1.error[ 787] = 1'b0;frame1.data[ 788] = 8'h09; frame1.valid[ 788] = 1'b1; frame1.error[ 788] = 1'b0;frame1.data[ 789] = 8'h0A; frame1.valid[ 789] = 1'b1; frame1.error[ 789] = 1'b0;frame1.data[ 790] = 8'h0B; frame1.valid[ 790] = 1'b1; frame1.error[ 790] = 1'b0;frame1.data[ 791] = 8'h0C; frame1.valid[ 791] = 1'b1; frame1.error[ 791] = 1'b0;frame1.data[ 792] = 8'h0D; frame1.valid[ 792] = 1'b1; frame1.error[ 792] = 1'b0;frame1.data[ 793] = 8'h0E; frame1.valid[ 793] = 1'b1; frame1.error[ 793] = 1'b0;frame1.data[ 794] = 8'h0F; frame1.valid[ 794] = 1'b1; frame1.error[ 794] = 1'b0;frame1.data[ 795] = 8'h10; frame1.valid[ 795] = 1'b1; frame1.error[ 795] = 1'b0;frame1.data[ 796] = 8'h11; frame1.valid[ 796] = 1'b1; frame1.error[ 796] = 1'b0;frame1.data[ 797] = 8'h12; frame1.valid[ 797] = 1'b1; frame1.error[ 797] = 1'b0;
        frame1.data[ 798] = 8'h13; frame1.valid[ 798] = 1'b1; frame1.error[ 798] = 1'b0;frame1.data[ 799] = 8'h14; frame1.valid[ 799] = 1'b1; frame1.error[ 799] = 1'b0;frame1.data[ 800] = 8'h15; frame1.valid[ 800] = 1'b1; frame1.error[ 800] = 1'b0;frame1.data[ 801] = 8'h16; frame1.valid[ 801] = 1'b1; frame1.error[ 801] = 1'b0;frame1.data[ 802] = 8'h17; frame1.valid[ 802] = 1'b1; frame1.error[ 802] = 1'b0;frame1.data[ 803] = 8'h18; frame1.valid[ 803] = 1'b1; frame1.error[ 803] = 1'b0;frame1.data[ 804] = 8'h19; frame1.valid[ 804] = 1'b1; frame1.error[ 804] = 1'b0;frame1.data[ 805] = 8'h1A; frame1.valid[ 805] = 1'b1; frame1.error[ 805] = 1'b0;frame1.data[ 806] = 8'h1B; frame1.valid[ 806] = 1'b1; frame1.error[ 806] = 1'b0;frame1.data[ 807] = 8'h1C; frame1.valid[ 807] = 1'b1; frame1.error[ 807] = 1'b0;frame1.data[ 808] = 8'h1D; frame1.valid[ 808] = 1'b1; frame1.error[ 808] = 1'b0;frame1.data[ 809] = 8'h1E; frame1.valid[ 809] = 1'b1; frame1.error[ 809] = 1'b0;frame1.data[ 810] = 8'h1F; frame1.valid[ 810] = 1'b1; frame1.error[ 810] = 1'b0;frame1.data[ 811] = 8'h20; frame1.valid[ 811] = 1'b1; frame1.error[ 811] = 1'b0;frame1.data[ 812] = 8'h21; frame1.valid[ 812] = 1'b1; frame1.error[ 812] = 1'b0;frame1.data[ 813] = 8'h22; frame1.valid[ 813] = 1'b1; frame1.error[ 813] = 1'b0;
        frame1.data[ 814] = 8'h23; frame1.valid[ 814] = 1'b1; frame1.error[ 814] = 1'b0;frame1.data[ 815] = 8'h24; frame1.valid[ 815] = 1'b1; frame1.error[ 815] = 1'b0;frame1.data[ 816] = 8'h25; frame1.valid[ 816] = 1'b1; frame1.error[ 816] = 1'b0;frame1.data[ 817] = 8'h26; frame1.valid[ 817] = 1'b1; frame1.error[ 817] = 1'b0;frame1.data[ 818] = 8'h27; frame1.valid[ 818] = 1'b1; frame1.error[ 818] = 1'b0;frame1.data[ 819] = 8'h28; frame1.valid[ 819] = 1'b1; frame1.error[ 819] = 1'b0;frame1.data[ 820] = 8'h29; frame1.valid[ 820] = 1'b1; frame1.error[ 820] = 1'b0;frame1.data[ 821] = 8'h2A; frame1.valid[ 821] = 1'b1; frame1.error[ 821] = 1'b0;frame1.data[ 822] = 8'h2B; frame1.valid[ 822] = 1'b1; frame1.error[ 822] = 1'b0;frame1.data[ 823] = 8'h2C; frame1.valid[ 823] = 1'b1; frame1.error[ 823] = 1'b0;frame1.data[ 824] = 8'h2D; frame1.valid[ 824] = 1'b1; frame1.error[ 824] = 1'b0;frame1.data[ 825] = 8'h2E; frame1.valid[ 825] = 1'b1; frame1.error[ 825] = 1'b0;frame1.data[ 826] = 8'h2F; frame1.valid[ 826] = 1'b1; frame1.error[ 826] = 1'b0;frame1.data[ 827] = 8'h30; frame1.valid[ 827] = 1'b1; frame1.error[ 827] = 1'b0;frame1.data[ 828] = 8'h31; frame1.valid[ 828] = 1'b1; frame1.error[ 828] = 1'b0;frame1.data[ 829] = 8'h32; frame1.valid[ 829] = 1'b1; frame1.error[ 829] = 1'b0;
        frame1.data[ 830] = 8'h33; frame1.valid[ 830] = 1'b1; frame1.error[ 830] = 1'b0;frame1.data[ 831] = 8'h34; frame1.valid[ 831] = 1'b1; frame1.error[ 831] = 1'b0;frame1.data[ 832] = 8'h35; frame1.valid[ 832] = 1'b1; frame1.error[ 832] = 1'b0;frame1.data[ 833] = 8'h36; frame1.valid[ 833] = 1'b1; frame1.error[ 833] = 1'b0;frame1.data[ 834] = 8'h37; frame1.valid[ 834] = 1'b1; frame1.error[ 834] = 1'b0;frame1.data[ 835] = 8'h38; frame1.valid[ 835] = 1'b1; frame1.error[ 835] = 1'b0;frame1.data[ 836] = 8'h39; frame1.valid[ 836] = 1'b1; frame1.error[ 836] = 1'b0;frame1.data[ 837] = 8'h3A; frame1.valid[ 837] = 1'b1; frame1.error[ 837] = 1'b0;frame1.data[ 838] = 8'h3B; frame1.valid[ 838] = 1'b1; frame1.error[ 838] = 1'b0;frame1.data[ 839] = 8'h3C; frame1.valid[ 839] = 1'b1; frame1.error[ 839] = 1'b0;frame1.data[ 840] = 8'h3D; frame1.valid[ 840] = 1'b1; frame1.error[ 840] = 1'b0;frame1.data[ 841] = 8'h3E; frame1.valid[ 841] = 1'b1; frame1.error[ 841] = 1'b0;frame1.data[ 842] = 8'h3F; frame1.valid[ 842] = 1'b1; frame1.error[ 842] = 1'b0;frame1.data[ 843] = 8'h40; frame1.valid[ 843] = 1'b1; frame1.error[ 843] = 1'b0;frame1.data[ 844] = 8'h41; frame1.valid[ 844] = 1'b1; frame1.error[ 844] = 1'b0;frame1.data[ 845] = 8'h42; frame1.valid[ 845] = 1'b1; frame1.error[ 845] = 1'b0;
        frame1.data[ 846] = 8'h43; frame1.valid[ 846] = 1'b1; frame1.error[ 846] = 1'b0;frame1.data[ 847] = 8'h44; frame1.valid[ 847] = 1'b1; frame1.error[ 847] = 1'b0;frame1.data[ 848] = 8'h45; frame1.valid[ 848] = 1'b1; frame1.error[ 848] = 1'b0;frame1.data[ 849] = 8'h46; frame1.valid[ 849] = 1'b1; frame1.error[ 849] = 1'b0;frame1.data[ 850] = 8'h47; frame1.valid[ 850] = 1'b1; frame1.error[ 850] = 1'b0;frame1.data[ 851] = 8'h48; frame1.valid[ 851] = 1'b1; frame1.error[ 851] = 1'b0;frame1.data[ 852] = 8'h49; frame1.valid[ 852] = 1'b1; frame1.error[ 852] = 1'b0;frame1.data[ 853] = 8'h4A; frame1.valid[ 853] = 1'b1; frame1.error[ 853] = 1'b0;frame1.data[ 854] = 8'h4B; frame1.valid[ 854] = 1'b1; frame1.error[ 854] = 1'b0;frame1.data[ 855] = 8'h4C; frame1.valid[ 855] = 1'b1; frame1.error[ 855] = 1'b0;frame1.data[ 856] = 8'h4D; frame1.valid[ 856] = 1'b1; frame1.error[ 856] = 1'b0;frame1.data[ 857] = 8'h4E; frame1.valid[ 857] = 1'b1; frame1.error[ 857] = 1'b0;frame1.data[ 858] = 8'h4F; frame1.valid[ 858] = 1'b1; frame1.error[ 858] = 1'b0;frame1.data[ 859] = 8'h50; frame1.valid[ 859] = 1'b1; frame1.error[ 859] = 1'b0;frame1.data[ 860] = 8'h51; frame1.valid[ 860] = 1'b1; frame1.error[ 860] = 1'b0;frame1.data[ 861] = 8'h52; frame1.valid[ 861] = 1'b1; frame1.error[ 861] = 1'b0;
        frame1.data[ 862] = 8'h53; frame1.valid[ 862] = 1'b1; frame1.error[ 862] = 1'b0;frame1.data[ 863] = 8'h54; frame1.valid[ 863] = 1'b1; frame1.error[ 863] = 1'b0;frame1.data[ 864] = 8'h55; frame1.valid[ 864] = 1'b1; frame1.error[ 864] = 1'b0;frame1.data[ 865] = 8'h56; frame1.valid[ 865] = 1'b1; frame1.error[ 865] = 1'b0;frame1.data[ 866] = 8'h57; frame1.valid[ 866] = 1'b1; frame1.error[ 866] = 1'b0;frame1.data[ 867] = 8'h58; frame1.valid[ 867] = 1'b1; frame1.error[ 867] = 1'b0;frame1.data[ 868] = 8'h59; frame1.valid[ 868] = 1'b1; frame1.error[ 868] = 1'b0;frame1.data[ 869] = 8'h5A; frame1.valid[ 869] = 1'b1; frame1.error[ 869] = 1'b0;frame1.data[ 870] = 8'h5B; frame1.valid[ 870] = 1'b1; frame1.error[ 870] = 1'b0;frame1.data[ 871] = 8'h5C; frame1.valid[ 871] = 1'b1; frame1.error[ 871] = 1'b0;frame1.data[ 872] = 8'h5D; frame1.valid[ 872] = 1'b1; frame1.error[ 872] = 1'b0;frame1.data[ 873] = 8'h5E; frame1.valid[ 873] = 1'b1; frame1.error[ 873] = 1'b0;frame1.data[ 874] = 8'h5F; frame1.valid[ 874] = 1'b1; frame1.error[ 874] = 1'b0;frame1.data[ 875] = 8'h60; frame1.valid[ 875] = 1'b1; frame1.error[ 875] = 1'b0;frame1.data[ 876] = 8'h61; frame1.valid[ 876] = 1'b1; frame1.error[ 876] = 1'b0;frame1.data[ 877] = 8'h62; frame1.valid[ 877] = 1'b1; frame1.error[ 877] = 1'b0;
        frame1.data[ 878] = 8'h63; frame1.valid[ 878] = 1'b1; frame1.error[ 878] = 1'b0;frame1.data[ 879] = 8'h64; frame1.valid[ 879] = 1'b1; frame1.error[ 879] = 1'b0;frame1.data[ 880] = 8'h65; frame1.valid[ 880] = 1'b1; frame1.error[ 880] = 1'b0;frame1.data[ 881] = 8'h66; frame1.valid[ 881] = 1'b1; frame1.error[ 881] = 1'b0;frame1.data[ 882] = 8'h67; frame1.valid[ 882] = 1'b1; frame1.error[ 882] = 1'b0;frame1.data[ 883] = 8'h68; frame1.valid[ 883] = 1'b1; frame1.error[ 883] = 1'b0;frame1.data[ 884] = 8'h69; frame1.valid[ 884] = 1'b1; frame1.error[ 884] = 1'b0;frame1.data[ 885] = 8'h6A; frame1.valid[ 885] = 1'b1; frame1.error[ 885] = 1'b0;frame1.data[ 886] = 8'h6B; frame1.valid[ 886] = 1'b1; frame1.error[ 886] = 1'b0;frame1.data[ 887] = 8'h6C; frame1.valid[ 887] = 1'b1; frame1.error[ 887] = 1'b0;frame1.data[ 888] = 8'h6D; frame1.valid[ 888] = 1'b1; frame1.error[ 888] = 1'b0;frame1.data[ 889] = 8'h6E; frame1.valid[ 889] = 1'b1; frame1.error[ 889] = 1'b0;frame1.data[ 890] = 8'h6F; frame1.valid[ 890] = 1'b1; frame1.error[ 890] = 1'b0;frame1.data[ 891] = 8'h70; frame1.valid[ 891] = 1'b1; frame1.error[ 891] = 1'b0;frame1.data[ 892] = 8'h71; frame1.valid[ 892] = 1'b1; frame1.error[ 892] = 1'b0;frame1.data[ 893] = 8'h72; frame1.valid[ 893] = 1'b1; frame1.error[ 893] = 1'b0;
        frame1.data[ 894] = 8'h73; frame1.valid[ 894] = 1'b1; frame1.error[ 894] = 1'b0;frame1.data[ 895] = 8'h74; frame1.valid[ 895] = 1'b1; frame1.error[ 895] = 1'b0;frame1.data[ 896] = 8'h75; frame1.valid[ 896] = 1'b1; frame1.error[ 896] = 1'b0;frame1.data[ 897] = 8'h76; frame1.valid[ 897] = 1'b1; frame1.error[ 897] = 1'b0;frame1.data[ 898] = 8'h77; frame1.valid[ 898] = 1'b1; frame1.error[ 898] = 1'b0;frame1.data[ 899] = 8'h78; frame1.valid[ 899] = 1'b1; frame1.error[ 899] = 1'b0;frame1.data[ 900] = 8'h79; frame1.valid[ 900] = 1'b1; frame1.error[ 900] = 1'b0;frame1.data[ 901] = 8'h7A; frame1.valid[ 901] = 1'b1; frame1.error[ 901] = 1'b0;frame1.data[ 902] = 8'h7B; frame1.valid[ 902] = 1'b1; frame1.error[ 902] = 1'b0;frame1.data[ 903] = 8'h7C; frame1.valid[ 903] = 1'b1; frame1.error[ 903] = 1'b0;frame1.data[ 904] = 8'h7D; frame1.valid[ 904] = 1'b1; frame1.error[ 904] = 1'b0;frame1.data[ 905] = 8'h7E; frame1.valid[ 905] = 1'b1; frame1.error[ 905] = 1'b0;frame1.data[ 906] = 8'h7F; frame1.valid[ 906] = 1'b1; frame1.error[ 906] = 1'b0;frame1.data[ 907] = 8'h80; frame1.valid[ 907] = 1'b1; frame1.error[ 907] = 1'b0;frame1.data[ 908] = 8'h81; frame1.valid[ 908] = 1'b1; frame1.error[ 908] = 1'b0;frame1.data[ 909] = 8'h82; frame1.valid[ 909] = 1'b1; frame1.error[ 909] = 1'b0;
        frame1.data[ 910] = 8'h83; frame1.valid[ 910] = 1'b1; frame1.error[ 910] = 1'b0;frame1.data[ 911] = 8'h84; frame1.valid[ 911] = 1'b1; frame1.error[ 911] = 1'b0;frame1.data[ 912] = 8'h85; frame1.valid[ 912] = 1'b1; frame1.error[ 912] = 1'b0;frame1.data[ 913] = 8'h86; frame1.valid[ 913] = 1'b1; frame1.error[ 913] = 1'b0;frame1.data[ 914] = 8'h87; frame1.valid[ 914] = 1'b1; frame1.error[ 914] = 1'b0;frame1.data[ 915] = 8'h88; frame1.valid[ 915] = 1'b1; frame1.error[ 915] = 1'b0;frame1.data[ 916] = 8'h89; frame1.valid[ 916] = 1'b1; frame1.error[ 916] = 1'b0;frame1.data[ 917] = 8'h8A; frame1.valid[ 917] = 1'b1; frame1.error[ 917] = 1'b0;frame1.data[ 918] = 8'h8B; frame1.valid[ 918] = 1'b1; frame1.error[ 918] = 1'b0;frame1.data[ 919] = 8'h8C; frame1.valid[ 919] = 1'b1; frame1.error[ 919] = 1'b0;frame1.data[ 920] = 8'h8D; frame1.valid[ 920] = 1'b1; frame1.error[ 920] = 1'b0;frame1.data[ 921] = 8'h8E; frame1.valid[ 921] = 1'b1; frame1.error[ 921] = 1'b0;frame1.data[ 922] = 8'h8F; frame1.valid[ 922] = 1'b1; frame1.error[ 922] = 1'b0;frame1.data[ 923] = 8'h90; frame1.valid[ 923] = 1'b1; frame1.error[ 923] = 1'b0;frame1.data[ 924] = 8'h91; frame1.valid[ 924] = 1'b1; frame1.error[ 924] = 1'b0;frame1.data[ 925] = 8'h92; frame1.valid[ 925] = 1'b1; frame1.error[ 925] = 1'b0;
        frame1.data[ 926] = 8'h93; frame1.valid[ 926] = 1'b1; frame1.error[ 926] = 1'b0;frame1.data[ 927] = 8'h94; frame1.valid[ 927] = 1'b1; frame1.error[ 927] = 1'b0;frame1.data[ 928] = 8'h95; frame1.valid[ 928] = 1'b1; frame1.error[ 928] = 1'b0;frame1.data[ 929] = 8'h96; frame1.valid[ 929] = 1'b1; frame1.error[ 929] = 1'b0;frame1.data[ 930] = 8'h97; frame1.valid[ 930] = 1'b1; frame1.error[ 930] = 1'b0;frame1.data[ 931] = 8'h98; frame1.valid[ 931] = 1'b1; frame1.error[ 931] = 1'b0;frame1.data[ 932] = 8'h99; frame1.valid[ 932] = 1'b1; frame1.error[ 932] = 1'b0;frame1.data[ 933] = 8'h9A; frame1.valid[ 933] = 1'b1; frame1.error[ 933] = 1'b0;frame1.data[ 934] = 8'h9B; frame1.valid[ 934] = 1'b1; frame1.error[ 934] = 1'b0;frame1.data[ 935] = 8'h9C; frame1.valid[ 935] = 1'b1; frame1.error[ 935] = 1'b0;frame1.data[ 936] = 8'h9D; frame1.valid[ 936] = 1'b1; frame1.error[ 936] = 1'b0;frame1.data[ 937] = 8'h9E; frame1.valid[ 937] = 1'b1; frame1.error[ 937] = 1'b0;frame1.data[ 938] = 8'h9F; frame1.valid[ 938] = 1'b1; frame1.error[ 938] = 1'b0;frame1.data[ 939] = 8'hA0; frame1.valid[ 939] = 1'b1; frame1.error[ 939] = 1'b0;frame1.data[ 940] = 8'hA1; frame1.valid[ 940] = 1'b1; frame1.error[ 940] = 1'b0;frame1.data[ 941] = 8'hA2; frame1.valid[ 941] = 1'b1; frame1.error[ 941] = 1'b0;
        frame1.data[ 942] = 8'hA3; frame1.valid[ 942] = 1'b1; frame1.error[ 942] = 1'b0;frame1.data[ 943] = 8'hA4; frame1.valid[ 943] = 1'b1; frame1.error[ 943] = 1'b0;frame1.data[ 944] = 8'hA5; frame1.valid[ 944] = 1'b1; frame1.error[ 944] = 1'b0;frame1.data[ 945] = 8'hA6; frame1.valid[ 945] = 1'b1; frame1.error[ 945] = 1'b0;frame1.data[ 946] = 8'hA7; frame1.valid[ 946] = 1'b1; frame1.error[ 946] = 1'b0;frame1.data[ 947] = 8'hA8; frame1.valid[ 947] = 1'b1; frame1.error[ 947] = 1'b0;frame1.data[ 948] = 8'hA9; frame1.valid[ 948] = 1'b1; frame1.error[ 948] = 1'b0;frame1.data[ 949] = 8'hAA; frame1.valid[ 949] = 1'b1; frame1.error[ 949] = 1'b0;frame1.data[ 950] = 8'hAB; frame1.valid[ 950] = 1'b1; frame1.error[ 950] = 1'b0;frame1.data[ 951] = 8'hAC; frame1.valid[ 951] = 1'b1; frame1.error[ 951] = 1'b0;frame1.data[ 952] = 8'hAD; frame1.valid[ 952] = 1'b1; frame1.error[ 952] = 1'b0;frame1.data[ 953] = 8'hAE; frame1.valid[ 953] = 1'b1; frame1.error[ 953] = 1'b0;frame1.data[ 954] = 8'hAF; frame1.valid[ 954] = 1'b1; frame1.error[ 954] = 1'b0;frame1.data[ 955] = 8'hB0; frame1.valid[ 955] = 1'b1; frame1.error[ 955] = 1'b0;frame1.data[ 956] = 8'hB1; frame1.valid[ 956] = 1'b1; frame1.error[ 956] = 1'b0;frame1.data[ 957] = 8'hB2; frame1.valid[ 957] = 1'b1; frame1.error[ 957] = 1'b0;
        frame1.data[ 958] = 8'hB3; frame1.valid[ 958] = 1'b1; frame1.error[ 958] = 1'b0;frame1.data[ 959] = 8'hB4; frame1.valid[ 959] = 1'b1; frame1.error[ 959] = 1'b0;frame1.data[ 960] = 8'hB5; frame1.valid[ 960] = 1'b1; frame1.error[ 960] = 1'b0;frame1.data[ 961] = 8'hB6; frame1.valid[ 961] = 1'b1; frame1.error[ 961] = 1'b0;frame1.data[ 962] = 8'hB7; frame1.valid[ 962] = 1'b1; frame1.error[ 962] = 1'b0;frame1.data[ 963] = 8'hB8; frame1.valid[ 963] = 1'b1; frame1.error[ 963] = 1'b0;frame1.data[ 964] = 8'hB9; frame1.valid[ 964] = 1'b1; frame1.error[ 964] = 1'b0;frame1.data[ 965] = 8'hBA; frame1.valid[ 965] = 1'b1; frame1.error[ 965] = 1'b0;frame1.data[ 966] = 8'hBB; frame1.valid[ 966] = 1'b1; frame1.error[ 966] = 1'b0;frame1.data[ 967] = 8'hBC; frame1.valid[ 967] = 1'b1; frame1.error[ 967] = 1'b0;frame1.data[ 968] = 8'hBD; frame1.valid[ 968] = 1'b1; frame1.error[ 968] = 1'b0;frame1.data[ 969] = 8'hBE; frame1.valid[ 969] = 1'b1; frame1.error[ 969] = 1'b0;frame1.data[ 970] = 8'hBF; frame1.valid[ 970] = 1'b1; frame1.error[ 970] = 1'b0;frame1.data[ 971] = 8'hC0; frame1.valid[ 971] = 1'b1; frame1.error[ 971] = 1'b0;frame1.data[ 972] = 8'hC1; frame1.valid[ 972] = 1'b1; frame1.error[ 972] = 1'b0;frame1.data[ 973] = 8'hC2; frame1.valid[ 973] = 1'b1; frame1.error[ 973] = 1'b0;
        frame1.data[ 974] = 8'hC3; frame1.valid[ 974] = 1'b1; frame1.error[ 974] = 1'b0;frame1.data[ 975] = 8'hC4; frame1.valid[ 975] = 1'b1; frame1.error[ 975] = 1'b0;frame1.data[ 976] = 8'hC5; frame1.valid[ 976] = 1'b1; frame1.error[ 976] = 1'b0;frame1.data[ 977] = 8'hC6; frame1.valid[ 977] = 1'b1; frame1.error[ 977] = 1'b0;frame1.data[ 978] = 8'hC7; frame1.valid[ 978] = 1'b1; frame1.error[ 978] = 1'b0;frame1.data[ 979] = 8'hC8; frame1.valid[ 979] = 1'b1; frame1.error[ 979] = 1'b0;frame1.data[ 980] = 8'hC9; frame1.valid[ 980] = 1'b1; frame1.error[ 980] = 1'b0;frame1.data[ 981] = 8'hCA; frame1.valid[ 981] = 1'b1; frame1.error[ 981] = 1'b0;frame1.data[ 982] = 8'hCB; frame1.valid[ 982] = 1'b1; frame1.error[ 982] = 1'b0;frame1.data[ 983] = 8'hCC; frame1.valid[ 983] = 1'b1; frame1.error[ 983] = 1'b0;frame1.data[ 984] = 8'hCD; frame1.valid[ 984] = 1'b1; frame1.error[ 984] = 1'b0;frame1.data[ 985] = 8'hCE; frame1.valid[ 985] = 1'b1; frame1.error[ 985] = 1'b0;frame1.data[ 986] = 8'hCF; frame1.valid[ 986] = 1'b1; frame1.error[ 986] = 1'b0;frame1.data[ 987] = 8'hD0; frame1.valid[ 987] = 1'b1; frame1.error[ 987] = 1'b0;frame1.data[ 988] = 8'hD1; frame1.valid[ 988] = 1'b1; frame1.error[ 988] = 1'b0;frame1.data[ 989] = 8'hD2; frame1.valid[ 989] = 1'b1; frame1.error[ 989] = 1'b0;
        frame1.data[ 990] = 8'hD3; frame1.valid[ 990] = 1'b1; frame1.error[ 990] = 1'b0;frame1.data[ 991] = 8'hD4; frame1.valid[ 991] = 1'b1; frame1.error[ 991] = 1'b0;frame1.data[ 992] = 8'hD5; frame1.valid[ 992] = 1'b1; frame1.error[ 992] = 1'b0;frame1.data[ 993] = 8'hD6; frame1.valid[ 993] = 1'b1; frame1.error[ 993] = 1'b0;frame1.data[ 994] = 8'hD7; frame1.valid[ 994] = 1'b1; frame1.error[ 994] = 1'b0;frame1.data[ 995] = 8'hD8; frame1.valid[ 995] = 1'b1; frame1.error[ 995] = 1'b0;frame1.data[ 996] = 8'hD9; frame1.valid[ 996] = 1'b1; frame1.error[ 996] = 1'b0;frame1.data[ 997] = 8'hDA; frame1.valid[ 997] = 1'b1; frame1.error[ 997] = 1'b0;frame1.data[ 998] = 8'hDB; frame1.valid[ 998] = 1'b1; frame1.error[ 998] = 1'b0;frame1.data[ 999] = 8'hDC; frame1.valid[ 999] = 1'b1; frame1.error[ 999] = 1'b0;frame1.data[1000] = 8'hDD; frame1.valid[1000] = 1'b1; frame1.error[1000] = 1'b0;frame1.data[1001] = 8'hDE; frame1.valid[1001] = 1'b1; frame1.error[1001] = 1'b0;frame1.data[1002] = 8'hDF; frame1.valid[1002] = 1'b1; frame1.error[1002] = 1'b0;frame1.data[1003] = 8'hE0; frame1.valid[1003] = 1'b1; frame1.error[1003] = 1'b0;frame1.data[1004] = 8'hE1; frame1.valid[1004] = 1'b1; frame1.error[1004] = 1'b0;frame1.data[1005] = 8'hE2; frame1.valid[1005] = 1'b1; frame1.error[1005] = 1'b0;
        frame1.data[1006] = 8'hE3; frame1.valid[1006] = 1'b1; frame1.error[1006] = 1'b0;frame1.data[1007] = 8'hE4; frame1.valid[1007] = 1'b1; frame1.error[1007] = 1'b0;frame1.data[1008] = 8'hE5; frame1.valid[1008] = 1'b1; frame1.error[1008] = 1'b0;frame1.data[1009] = 8'hE6; frame1.valid[1009] = 1'b1; frame1.error[1009] = 1'b0;frame1.data[1010] = 8'hE7; frame1.valid[1010] = 1'b1; frame1.error[1010] = 1'b0;frame1.data[1011] = 8'hE8; frame1.valid[1011] = 1'b1; frame1.error[1011] = 1'b0;frame1.data[1012] = 8'hE9; frame1.valid[1012] = 1'b1; frame1.error[1012] = 1'b0;frame1.data[1013] = 8'hEA; frame1.valid[1013] = 1'b1; frame1.error[1013] = 1'b0;frame1.data[1014] = 8'hEB; frame1.valid[1014] = 1'b1; frame1.error[1014] = 1'b0;frame1.data[1015] = 8'hEC; frame1.valid[1015] = 1'b1; frame1.error[1015] = 1'b0;frame1.data[1016] = 8'hED; frame1.valid[1016] = 1'b1; frame1.error[1016] = 1'b0;frame1.data[1017] = 8'hEE; frame1.valid[1017] = 1'b1; frame1.error[1017] = 1'b0;frame1.data[1018] = 8'hEF; frame1.valid[1018] = 1'b1; frame1.error[1018] = 1'b0;frame1.data[1019] = 8'hF0; frame1.valid[1019] = 1'b1; frame1.error[1019] = 1'b0;frame1.data[1020] = 8'hF1; frame1.valid[1020] = 1'b1; frame1.error[1020] = 1'b0;frame1.data[1021] = 8'hF2; frame1.valid[1021] = 1'b1; frame1.error[1021] = 1'b0;
        frame1.data[1022] = 8'hF3; frame1.valid[1022] = 1'b1; frame1.error[1022] = 1'b0;frame1.data[1023] = 8'hF4; frame1.valid[1023] = 1'b1; frame1.error[1023] = 1'b0;frame1.data[1024] = 8'hF5; frame1.valid[1024] = 1'b1; frame1.error[1024] = 1'b0;frame1.data[1025] = 8'hF6; frame1.valid[1025] = 1'b1; frame1.error[1025] = 1'b0;frame1.data[1026] = 8'hF7; frame1.valid[1026] = 1'b1; frame1.error[1026] = 1'b0;frame1.data[1027] = 8'hF8; frame1.valid[1027] = 1'b1; frame1.error[1027] = 1'b0;frame1.data[1028] = 8'hF9; frame1.valid[1028] = 1'b1; frame1.error[1028] = 1'b0;frame1.data[1029] = 8'hFA; frame1.valid[1029] = 1'b1; frame1.error[1029] = 1'b0;frame1.data[1030] = 8'hFB; frame1.valid[1030] = 1'b1; frame1.error[1030] = 1'b0;frame1.data[1031] = 8'hFC; frame1.valid[1031] = 1'b1; frame1.error[1031] = 1'b0;frame1.data[1032] = 8'hFD; frame1.valid[1032] = 1'b1; frame1.error[1032] = 1'b0;frame1.data[1033] = 8'hFE; frame1.valid[1033] = 1'b1; frame1.error[1033] = 1'b0;frame1.data[1034] = 8'h00; frame1.valid[1034] = 1'b1; frame1.error[1034] = 1'b0;frame1.data[1035] = 8'h01; frame1.valid[1035] = 1'b1; frame1.error[1035] = 1'b0;frame1.data[1036] = 8'h02; frame1.valid[1036] = 1'b1; frame1.error[1036] = 1'b0;frame1.data[1037] = 8'h03; frame1.valid[1037] = 1'b1; frame1.error[1037] = 1'b0;
        frame1.data[1038] = 8'h04; frame1.valid[1038] = 1'b1; frame1.error[1038] = 1'b0;frame1.data[1039] = 8'h05; frame1.valid[1039] = 1'b1; frame1.error[1039] = 1'b0;frame1.data[1040] = 8'h06; frame1.valid[1040] = 1'b1; frame1.error[1040] = 1'b0;frame1.data[1041] = 8'h07; frame1.valid[1041] = 1'b1; frame1.error[1041] = 1'b0;frame1.data[1042] = 8'h08; frame1.valid[1042] = 1'b1; frame1.error[1042] = 1'b0;frame1.data[1043] = 8'h09; frame1.valid[1043] = 1'b1; frame1.error[1043] = 1'b0;frame1.data[1044] = 8'h0A; frame1.valid[1044] = 1'b1; frame1.error[1044] = 1'b0;frame1.data[1045] = 8'h0B; frame1.valid[1045] = 1'b1; frame1.error[1045] = 1'b0;frame1.data[1046] = 8'h0C; frame1.valid[1046] = 1'b1; frame1.error[1046] = 1'b0;frame1.data[1047] = 8'h0D; frame1.valid[1047] = 1'b1; frame1.error[1047] = 1'b0;frame1.data[1048] = 8'h0E; frame1.valid[1048] = 1'b1; frame1.error[1048] = 1'b0;frame1.data[1049] = 8'h0F; frame1.valid[1049] = 1'b1; frame1.error[1049] = 1'b0;frame1.data[1050] = 8'h10; frame1.valid[1050] = 1'b1; frame1.error[1050] = 1'b0;frame1.data[1051] = 8'h11; frame1.valid[1051] = 1'b1; frame1.error[1051] = 1'b0;frame1.data[1052] = 8'h12; frame1.valid[1052] = 1'b1; frame1.error[1052] = 1'b0;frame1.data[1053] = 8'h13; frame1.valid[1053] = 1'b1; frame1.error[1053] = 1'b0;
        frame1.data[1054] = 8'h14; frame1.valid[1054] = 1'b1; frame1.error[1054] = 1'b0;frame1.data[1055] = 8'h15; frame1.valid[1055] = 1'b1; frame1.error[1055] = 1'b0;frame1.data[1056] = 8'h16; frame1.valid[1056] = 1'b1; frame1.error[1056] = 1'b0;frame1.data[1057] = 8'h17; frame1.valid[1057] = 1'b1; frame1.error[1057] = 1'b0;frame1.data[1058] = 8'h18; frame1.valid[1058] = 1'b1; frame1.error[1058] = 1'b0;frame1.data[1059] = 8'h19; frame1.valid[1059] = 1'b1; frame1.error[1059] = 1'b0;frame1.data[1060] = 8'h1A; frame1.valid[1060] = 1'b1; frame1.error[1060] = 1'b0;frame1.data[1061] = 8'h1B; frame1.valid[1061] = 1'b1; frame1.error[1061] = 1'b0;frame1.data[1062] = 8'h1C; frame1.valid[1062] = 1'b1; frame1.error[1062] = 1'b0;frame1.data[1063] = 8'h1D; frame1.valid[1063] = 1'b1; frame1.error[1063] = 1'b0;frame1.data[1064] = 8'h1E; frame1.valid[1064] = 1'b1; frame1.error[1064] = 1'b0;frame1.data[1065] = 8'h1F; frame1.valid[1065] = 1'b1; frame1.error[1065] = 1'b0;frame1.data[1066] = 8'h20; frame1.valid[1066] = 1'b1; frame1.error[1066] = 1'b0;frame1.data[1067] = 8'h21; frame1.valid[1067] = 1'b1; frame1.error[1067] = 1'b0;frame1.data[1068] = 8'h22; frame1.valid[1068] = 1'b1; frame1.error[1068] = 1'b0;frame1.data[1069] = 8'h23; frame1.valid[1069] = 1'b1; frame1.error[1069] = 1'b0;
        frame1.data[1070] = 8'h24; frame1.valid[1070] = 1'b1; frame1.error[1070] = 1'b0;frame1.data[1071] = 8'h25; frame1.valid[1071] = 1'b1; frame1.error[1071] = 1'b0;frame1.data[1072] = 8'h26; frame1.valid[1072] = 1'b1; frame1.error[1072] = 1'b0;frame1.data[1073] = 8'h27; frame1.valid[1073] = 1'b1; frame1.error[1073] = 1'b0;frame1.data[1074] = 8'h28; frame1.valid[1074] = 1'b1; frame1.error[1074] = 1'b0;frame1.data[1075] = 8'h29; frame1.valid[1075] = 1'b1; frame1.error[1075] = 1'b0;frame1.data[1076] = 8'h2A; frame1.valid[1076] = 1'b1; frame1.error[1076] = 1'b0;frame1.data[1077] = 8'h2B; frame1.valid[1077] = 1'b1; frame1.error[1077] = 1'b0;frame1.data[1078] = 8'h2C; frame1.valid[1078] = 1'b1; frame1.error[1078] = 1'b0;frame1.data[1079] = 8'h2D; frame1.valid[1079] = 1'b1; frame1.error[1079] = 1'b0;frame1.data[1080] = 8'h2E; frame1.valid[1080] = 1'b1; frame1.error[1080] = 1'b0;frame1.data[1081] = 8'h2F; frame1.valid[1081] = 1'b1; frame1.error[1081] = 1'b0;frame1.data[1082] = 8'h30; frame1.valid[1082] = 1'b1; frame1.error[1082] = 1'b0;frame1.data[1083] = 8'h31; frame1.valid[1083] = 1'b1; frame1.error[1083] = 1'b0;frame1.data[1084] = 8'h32; frame1.valid[1084] = 1'b1; frame1.error[1084] = 1'b0;frame1.data[1085] = 8'h33; frame1.valid[1085] = 1'b1; frame1.error[1085] = 1'b0;
        frame1.data[1086] = 8'h34; frame1.valid[1086] = 1'b1; frame1.error[1086] = 1'b0;frame1.data[1087] = 8'h35; frame1.valid[1087] = 1'b1; frame1.error[1087] = 1'b0;frame1.data[1088] = 8'h36; frame1.valid[1088] = 1'b1; frame1.error[1088] = 1'b0;frame1.data[1089] = 8'h37; frame1.valid[1089] = 1'b1; frame1.error[1089] = 1'b0;frame1.data[1090] = 8'h38; frame1.valid[1090] = 1'b1; frame1.error[1090] = 1'b0;frame1.data[1091] = 8'h39; frame1.valid[1091] = 1'b1; frame1.error[1091] = 1'b0;frame1.data[1092] = 8'h3A; frame1.valid[1092] = 1'b1; frame1.error[1092] = 1'b0;frame1.data[1093] = 8'h3B; frame1.valid[1093] = 1'b1; frame1.error[1093] = 1'b0;frame1.data[1094] = 8'h3C; frame1.valid[1094] = 1'b1; frame1.error[1094] = 1'b0;frame1.data[1095] = 8'h3D; frame1.valid[1095] = 1'b1; frame1.error[1095] = 1'b0;frame1.data[1096] = 8'h3E; frame1.valid[1096] = 1'b1; frame1.error[1096] = 1'b0;frame1.data[1097] = 8'h3F; frame1.valid[1097] = 1'b1; frame1.error[1097] = 1'b0;frame1.data[1098] = 8'h40; frame1.valid[1098] = 1'b1; frame1.error[1098] = 1'b0;frame1.data[1099] = 8'h41; frame1.valid[1099] = 1'b1; frame1.error[1099] = 1'b0;frame1.data[1100] = 8'h42; frame1.valid[1100] = 1'b1; frame1.error[1100] = 1'b0;frame1.data[1101] = 8'h43; frame1.valid[1101] = 1'b1; frame1.error[1101] = 1'b0;
        frame1.data[1102] = 8'h44; frame1.valid[1102] = 1'b1; frame1.error[1102] = 1'b0;frame1.data[1103] = 8'h45; frame1.valid[1103] = 1'b1; frame1.error[1103] = 1'b0;frame1.data[1104] = 8'h46; frame1.valid[1104] = 1'b1; frame1.error[1104] = 1'b0;frame1.data[1105] = 8'h47; frame1.valid[1105] = 1'b1; frame1.error[1105] = 1'b0;frame1.data[1106] = 8'h48; frame1.valid[1106] = 1'b1; frame1.error[1106] = 1'b0;frame1.data[1107] = 8'h49; frame1.valid[1107] = 1'b1; frame1.error[1107] = 1'b0;frame1.data[1108] = 8'h4A; frame1.valid[1108] = 1'b1; frame1.error[1108] = 1'b0;frame1.data[1109] = 8'h4B; frame1.valid[1109] = 1'b1; frame1.error[1109] = 1'b0;frame1.data[1110] = 8'h4C; frame1.valid[1110] = 1'b1; frame1.error[1110] = 1'b0;frame1.data[1111] = 8'h4D; frame1.valid[1111] = 1'b1; frame1.error[1111] = 1'b0;frame1.data[1112] = 8'h4E; frame1.valid[1112] = 1'b1; frame1.error[1112] = 1'b0;frame1.data[1113] = 8'h4F; frame1.valid[1113] = 1'b1; frame1.error[1113] = 1'b0;frame1.data[1114] = 8'h50; frame1.valid[1114] = 1'b1; frame1.error[1114] = 1'b0;frame1.data[1115] = 8'h51; frame1.valid[1115] = 1'b1; frame1.error[1115] = 1'b0;frame1.data[1116] = 8'h52; frame1.valid[1116] = 1'b1; frame1.error[1116] = 1'b0;frame1.data[1117] = 8'h53; frame1.valid[1117] = 1'b1; frame1.error[1117] = 1'b0;
        frame1.data[1118] = 8'h54; frame1.valid[1118] = 1'b1; frame1.error[1118] = 1'b0;frame1.data[1119] = 8'h55; frame1.valid[1119] = 1'b1; frame1.error[1119] = 1'b0;frame1.data[1120] = 8'h56; frame1.valid[1120] = 1'b1; frame1.error[1120] = 1'b0;frame1.data[1121] = 8'h57; frame1.valid[1121] = 1'b1; frame1.error[1121] = 1'b0;frame1.data[1122] = 8'h58; frame1.valid[1122] = 1'b1; frame1.error[1122] = 1'b0;frame1.data[1123] = 8'h59; frame1.valid[1123] = 1'b1; frame1.error[1123] = 1'b0;frame1.data[1124] = 8'h5A; frame1.valid[1124] = 1'b1; frame1.error[1124] = 1'b0;frame1.data[1125] = 8'h5B; frame1.valid[1125] = 1'b1; frame1.error[1125] = 1'b0;frame1.data[1126] = 8'h5C; frame1.valid[1126] = 1'b1; frame1.error[1126] = 1'b0;frame1.data[1127] = 8'h5D; frame1.valid[1127] = 1'b1; frame1.error[1127] = 1'b0;frame1.data[1128] = 8'h5E; frame1.valid[1128] = 1'b1; frame1.error[1128] = 1'b0;frame1.data[1129] = 8'h5F; frame1.valid[1129] = 1'b1; frame1.error[1129] = 1'b0;frame1.data[1130] = 8'h60; frame1.valid[1130] = 1'b1; frame1.error[1130] = 1'b0;frame1.data[1131] = 8'h61; frame1.valid[1131] = 1'b1; frame1.error[1131] = 1'b0;frame1.data[1132] = 8'h62; frame1.valid[1132] = 1'b1; frame1.error[1132] = 1'b0;frame1.data[1133] = 8'h63; frame1.valid[1133] = 1'b1; frame1.error[1133] = 1'b0;
        frame1.data[1134] = 8'h64; frame1.valid[1134] = 1'b1; frame1.error[1134] = 1'b0;frame1.data[1135] = 8'h65; frame1.valid[1135] = 1'b1; frame1.error[1135] = 1'b0;frame1.data[1136] = 8'h66; frame1.valid[1136] = 1'b1; frame1.error[1136] = 1'b0;frame1.data[1137] = 8'h67; frame1.valid[1137] = 1'b1; frame1.error[1137] = 1'b0;frame1.data[1138] = 8'h68; frame1.valid[1138] = 1'b1; frame1.error[1138] = 1'b0;frame1.data[1139] = 8'h69; frame1.valid[1139] = 1'b1; frame1.error[1139] = 1'b0;frame1.data[1140] = 8'h6A; frame1.valid[1140] = 1'b1; frame1.error[1140] = 1'b0;frame1.data[1141] = 8'h6B; frame1.valid[1141] = 1'b1; frame1.error[1141] = 1'b0;frame1.data[1142] = 8'h6C; frame1.valid[1142] = 1'b1; frame1.error[1142] = 1'b0;frame1.data[1143] = 8'h6D; frame1.valid[1143] = 1'b1; frame1.error[1143] = 1'b0;frame1.data[1144] = 8'h6E; frame1.valid[1144] = 1'b1; frame1.error[1144] = 1'b0;frame1.data[1145] = 8'h6F; frame1.valid[1145] = 1'b1; frame1.error[1145] = 1'b0;frame1.data[1146] = 8'h70; frame1.valid[1146] = 1'b1; frame1.error[1146] = 1'b0;frame1.data[1147] = 8'h71; frame1.valid[1147] = 1'b1; frame1.error[1147] = 1'b0;frame1.data[1148] = 8'h72; frame1.valid[1148] = 1'b1; frame1.error[1148] = 1'b0;frame1.data[1149] = 8'h73; frame1.valid[1149] = 1'b1; frame1.error[1149] = 1'b0;
        frame1.data[1150] = 8'h74; frame1.valid[1150] = 1'b1; frame1.error[1150] = 1'b0;frame1.data[1151] = 8'h75; frame1.valid[1151] = 1'b1; frame1.error[1151] = 1'b0;frame1.data[1152] = 8'h76; frame1.valid[1152] = 1'b1; frame1.error[1152] = 1'b0;frame1.data[1153] = 8'h77; frame1.valid[1153] = 1'b1; frame1.error[1153] = 1'b0;frame1.data[1154] = 8'h78; frame1.valid[1154] = 1'b1; frame1.error[1154] = 1'b0;frame1.data[1155] = 8'h79; frame1.valid[1155] = 1'b1; frame1.error[1155] = 1'b0;frame1.data[1156] = 8'h7A; frame1.valid[1156] = 1'b1; frame1.error[1156] = 1'b0;frame1.data[1157] = 8'h7B; frame1.valid[1157] = 1'b1; frame1.error[1157] = 1'b0;frame1.data[1158] = 8'h7C; frame1.valid[1158] = 1'b1; frame1.error[1158] = 1'b0;frame1.data[1159] = 8'h7D; frame1.valid[1159] = 1'b1; frame1.error[1159] = 1'b0;frame1.data[1160] = 8'h7E; frame1.valid[1160] = 1'b1; frame1.error[1160] = 1'b0;frame1.data[1161] = 8'h7F; frame1.valid[1161] = 1'b1; frame1.error[1161] = 1'b0;frame1.data[1162] = 8'h80; frame1.valid[1162] = 1'b1; frame1.error[1162] = 1'b0;frame1.data[1163] = 8'h81; frame1.valid[1163] = 1'b1; frame1.error[1163] = 1'b0;frame1.data[1164] = 8'h82; frame1.valid[1164] = 1'b1; frame1.error[1164] = 1'b0;frame1.data[1165] = 8'h83; frame1.valid[1165] = 1'b1; frame1.error[1165] = 1'b0;
        frame1.data[1166] = 8'h84; frame1.valid[1166] = 1'b1; frame1.error[1166] = 1'b0;frame1.data[1167] = 8'h85; frame1.valid[1167] = 1'b1; frame1.error[1167] = 1'b0;frame1.data[1168] = 8'h86; frame1.valid[1168] = 1'b1; frame1.error[1168] = 1'b0;frame1.data[1169] = 8'h87; frame1.valid[1169] = 1'b1; frame1.error[1169] = 1'b0;frame1.data[1170] = 8'h88; frame1.valid[1170] = 1'b1; frame1.error[1170] = 1'b0;frame1.data[1171] = 8'h89; frame1.valid[1171] = 1'b1; frame1.error[1171] = 1'b0;frame1.data[1172] = 8'h8A; frame1.valid[1172] = 1'b1; frame1.error[1172] = 1'b0;frame1.data[1173] = 8'h8B; frame1.valid[1173] = 1'b1; frame1.error[1173] = 1'b0;frame1.data[1174] = 8'h8C; frame1.valid[1174] = 1'b1; frame1.error[1174] = 1'b0;frame1.data[1175] = 8'h8D; frame1.valid[1175] = 1'b1; frame1.error[1175] = 1'b0;frame1.data[1176] = 8'h8E; frame1.valid[1176] = 1'b1; frame1.error[1176] = 1'b0;frame1.data[1177] = 8'h8F; frame1.valid[1177] = 1'b1; frame1.error[1177] = 1'b0;frame1.data[1178] = 8'h90; frame1.valid[1178] = 1'b1; frame1.error[1178] = 1'b0;frame1.data[1179] = 8'h91; frame1.valid[1179] = 1'b1; frame1.error[1179] = 1'b0;frame1.data[1180] = 8'h92; frame1.valid[1180] = 1'b1; frame1.error[1180] = 1'b0;frame1.data[1181] = 8'h93; frame1.valid[1181] = 1'b1; frame1.error[1181] = 1'b0;
        frame1.data[1182] = 8'h94; frame1.valid[1182] = 1'b1; frame1.error[1182] = 1'b0;frame1.data[1183] = 8'h95; frame1.valid[1183] = 1'b1; frame1.error[1183] = 1'b0;frame1.data[1184] = 8'h96; frame1.valid[1184] = 1'b1; frame1.error[1184] = 1'b0;frame1.data[1185] = 8'h97; frame1.valid[1185] = 1'b1; frame1.error[1185] = 1'b0;frame1.data[1186] = 8'h98; frame1.valid[1186] = 1'b1; frame1.error[1186] = 1'b0;frame1.data[1187] = 8'h99; frame1.valid[1187] = 1'b1; frame1.error[1187] = 1'b0;frame1.data[1188] = 8'h9A; frame1.valid[1188] = 1'b1; frame1.error[1188] = 1'b0;frame1.data[1189] = 8'h9B; frame1.valid[1189] = 1'b1; frame1.error[1189] = 1'b0;frame1.data[1190] = 8'h9C; frame1.valid[1190] = 1'b1; frame1.error[1190] = 1'b0;frame1.data[1191] = 8'h9D; frame1.valid[1191] = 1'b1; frame1.error[1191] = 1'b0;frame1.data[1192] = 8'h9E; frame1.valid[1192] = 1'b1; frame1.error[1192] = 1'b0;frame1.data[1193] = 8'h9F; frame1.valid[1193] = 1'b1; frame1.error[1193] = 1'b0;frame1.data[1194] = 8'hA0; frame1.valid[1194] = 1'b1; frame1.error[1194] = 1'b0;frame1.data[1195] = 8'hA1; frame1.valid[1195] = 1'b1; frame1.error[1195] = 1'b0;frame1.data[1196] = 8'hA2; frame1.valid[1196] = 1'b1; frame1.error[1196] = 1'b0;frame1.data[1197] = 8'hA3; frame1.valid[1197] = 1'b1; frame1.error[1197] = 1'b0;
        frame1.data[1198] = 8'hA4; frame1.valid[1198] = 1'b1; frame1.error[1198] = 1'b0;frame1.data[1199] = 8'hA5; frame1.valid[1199] = 1'b1; frame1.error[1199] = 1'b0;frame1.data[1200] = 8'hA6; frame1.valid[1200] = 1'b1; frame1.error[1200] = 1'b0;frame1.data[1201] = 8'hA7; frame1.valid[1201] = 1'b1; frame1.error[1201] = 1'b0;frame1.data[1202] = 8'hA8; frame1.valid[1202] = 1'b1; frame1.error[1202] = 1'b0;frame1.data[1203] = 8'hA9; frame1.valid[1203] = 1'b1; frame1.error[1203] = 1'b0;frame1.data[1204] = 8'hAA; frame1.valid[1204] = 1'b1; frame1.error[1204] = 1'b0;frame1.data[1205] = 8'hAB; frame1.valid[1205] = 1'b1; frame1.error[1205] = 1'b0;frame1.data[1206] = 8'hAC; frame1.valid[1206] = 1'b1; frame1.error[1206] = 1'b0;frame1.data[1207] = 8'hAD; frame1.valid[1207] = 1'b1; frame1.error[1207] = 1'b0;frame1.data[1208] = 8'hAE; frame1.valid[1208] = 1'b1; frame1.error[1208] = 1'b0;frame1.data[1209] = 8'hAF; frame1.valid[1209] = 1'b1; frame1.error[1209] = 1'b0;frame1.data[1210] = 8'hB0; frame1.valid[1210] = 1'b1; frame1.error[1210] = 1'b0;frame1.data[1211] = 8'hB1; frame1.valid[1211] = 1'b1; frame1.error[1211] = 1'b0;frame1.data[1212] = 8'hB2; frame1.valid[1212] = 1'b1; frame1.error[1212] = 1'b0;frame1.data[1213] = 8'hB3; frame1.valid[1213] = 1'b1; frame1.error[1213] = 1'b0;
        frame1.data[1214] = 8'hB4; frame1.valid[1214] = 1'b1; frame1.error[1214] = 1'b0;frame1.data[1215] = 8'hB5; frame1.valid[1215] = 1'b1; frame1.error[1215] = 1'b0;frame1.data[1216] = 8'hB6; frame1.valid[1216] = 1'b1; frame1.error[1216] = 1'b0;frame1.data[1217] = 8'hB7; frame1.valid[1217] = 1'b1; frame1.error[1217] = 1'b0;frame1.data[1218] = 8'hB8; frame1.valid[1218] = 1'b1; frame1.error[1218] = 1'b0;frame1.data[1219] = 8'hB9; frame1.valid[1219] = 1'b1; frame1.error[1219] = 1'b0;frame1.data[1220] = 8'hBA; frame1.valid[1220] = 1'b1; frame1.error[1220] = 1'b0;frame1.data[1221] = 8'hBB; frame1.valid[1221] = 1'b1; frame1.error[1221] = 1'b0;frame1.data[1222] = 8'hBC; frame1.valid[1222] = 1'b1; frame1.error[1222] = 1'b0;frame1.data[1223] = 8'hBD; frame1.valid[1223] = 1'b1; frame1.error[1223] = 1'b0;frame1.data[1224] = 8'hBE; frame1.valid[1224] = 1'b1; frame1.error[1224] = 1'b0;frame1.data[1225] = 8'hBF; frame1.valid[1225] = 1'b1; frame1.error[1225] = 1'b0;frame1.data[1226] = 8'hC0; frame1.valid[1226] = 1'b1; frame1.error[1226] = 1'b0;frame1.data[1227] = 8'hC1; frame1.valid[1227] = 1'b1; frame1.error[1227] = 1'b0;frame1.data[1228] = 8'hC2; frame1.valid[1228] = 1'b1; frame1.error[1228] = 1'b0;frame1.data[1229] = 8'hC3; frame1.valid[1229] = 1'b1; frame1.error[1229] = 1'b0;
        frame1.data[1230] = 8'hC4; frame1.valid[1230] = 1'b1; frame1.error[1230] = 1'b0;frame1.data[1231] = 8'hC5; frame1.valid[1231] = 1'b1; frame1.error[1231] = 1'b0;frame1.data[1232] = 8'hC6; frame1.valid[1232] = 1'b1; frame1.error[1232] = 1'b0;frame1.data[1233] = 8'hC7; frame1.valid[1233] = 1'b1; frame1.error[1233] = 1'b0;frame1.data[1234] = 8'hC8; frame1.valid[1234] = 1'b1; frame1.error[1234] = 1'b0;frame1.data[1235] = 8'hC9; frame1.valid[1235] = 1'b1; frame1.error[1235] = 1'b0;frame1.data[1236] = 8'hCA; frame1.valid[1236] = 1'b1; frame1.error[1236] = 1'b0;frame1.data[1237] = 8'hCB; frame1.valid[1237] = 1'b1; frame1.error[1237] = 1'b0;frame1.data[1238] = 8'hCC; frame1.valid[1238] = 1'b1; frame1.error[1238] = 1'b0;frame1.data[1239] = 8'hCD; frame1.valid[1239] = 1'b1; frame1.error[1239] = 1'b0;frame1.data[1240] = 8'hCE; frame1.valid[1240] = 1'b1; frame1.error[1240] = 1'b0;frame1.data[1241] = 8'hCF; frame1.valid[1241] = 1'b1; frame1.error[1241] = 1'b0;frame1.data[1242] = 8'hD0; frame1.valid[1242] = 1'b1; frame1.error[1242] = 1'b0;frame1.data[1243] = 8'hD1; frame1.valid[1243] = 1'b1; frame1.error[1243] = 1'b0;frame1.data[1244] = 8'hD2; frame1.valid[1244] = 1'b1; frame1.error[1244] = 1'b0;frame1.data[1245] = 8'hD3; frame1.valid[1245] = 1'b1; frame1.error[1245] = 1'b0;
        frame1.data[1246] = 8'hD4; frame1.valid[1246] = 1'b1; frame1.error[1246] = 1'b0;frame1.data[1247] = 8'hD5; frame1.valid[1247] = 1'b1; frame1.error[1247] = 1'b0;frame1.data[1248] = 8'hD6; frame1.valid[1248] = 1'b1; frame1.error[1248] = 1'b0;frame1.data[1249] = 8'hD7; frame1.valid[1249] = 1'b1; frame1.error[1249] = 1'b0;frame1.data[1250] = 8'hD8; frame1.valid[1250] = 1'b1; frame1.error[1250] = 1'b0;frame1.data[1251] = 8'hD9; frame1.valid[1251] = 1'b1; frame1.error[1251] = 1'b0;frame1.data[1252] = 8'hDA; frame1.valid[1252] = 1'b1; frame1.error[1252] = 1'b0;frame1.data[1253] = 8'hDB; frame1.valid[1253] = 1'b1; frame1.error[1253] = 1'b0;frame1.data[1254] = 8'hDC; frame1.valid[1254] = 1'b1; frame1.error[1254] = 1'b0;frame1.data[1255] = 8'hDD; frame1.valid[1255] = 1'b1; frame1.error[1255] = 1'b0;frame1.data[1256] = 8'hDE; frame1.valid[1256] = 1'b1; frame1.error[1256] = 1'b0;frame1.data[1257] = 8'hDF; frame1.valid[1257] = 1'b1; frame1.error[1257] = 1'b0;frame1.data[1258] = 8'hE0; frame1.valid[1258] = 1'b1; frame1.error[1258] = 1'b0;frame1.data[1259] = 8'hE1; frame1.valid[1259] = 1'b1; frame1.error[1259] = 1'b0;frame1.data[1260] = 8'hE2; frame1.valid[1260] = 1'b1; frame1.error[1260] = 1'b0;frame1.data[1261] = 8'hE3; frame1.valid[1261] = 1'b1; frame1.error[1261] = 1'b0;
        frame1.data[1262] = 8'hE4; frame1.valid[1262] = 1'b1; frame1.error[1262] = 1'b0;frame1.data[1263] = 8'hE5; frame1.valid[1263] = 1'b1; frame1.error[1263] = 1'b0;frame1.data[1264] = 8'hE6; frame1.valid[1264] = 1'b1; frame1.error[1264] = 1'b0;frame1.data[1265] = 8'hE7; frame1.valid[1265] = 1'b1; frame1.error[1265] = 1'b0;frame1.data[1266] = 8'hE8; frame1.valid[1266] = 1'b1; frame1.error[1266] = 1'b0;frame1.data[1267] = 8'hE9; frame1.valid[1267] = 1'b1; frame1.error[1267] = 1'b0;frame1.data[1268] = 8'hEA; frame1.valid[1268] = 1'b1; frame1.error[1268] = 1'b0;frame1.data[1269] = 8'hEB; frame1.valid[1269] = 1'b1; frame1.error[1269] = 1'b0;frame1.data[1270] = 8'hEC; frame1.valid[1270] = 1'b1; frame1.error[1270] = 1'b0;frame1.data[1271] = 8'hED; frame1.valid[1271] = 1'b1; frame1.error[1271] = 1'b0;frame1.data[1272] = 8'hEE; frame1.valid[1272] = 1'b1; frame1.error[1272] = 1'b0;frame1.data[1273] = 8'hEF; frame1.valid[1273] = 1'b1; frame1.error[1273] = 1'b0;frame1.data[1274] = 8'hF0; frame1.valid[1274] = 1'b1; frame1.error[1274] = 1'b0;frame1.data[1275] = 8'hF1; frame1.valid[1275] = 1'b1; frame1.error[1275] = 1'b0;frame1.data[1276] = 8'hF2; frame1.valid[1276] = 1'b1; frame1.error[1276] = 1'b0;frame1.data[1277] = 8'hF3; frame1.valid[1277] = 1'b1; frame1.error[1277] = 1'b0;
        frame1.data[1278] = 8'hF4; frame1.valid[1278] = 1'b1; frame1.error[1278] = 1'b0;frame1.data[1279] = 8'hF5; frame1.valid[1279] = 1'b1; frame1.error[1279] = 1'b0;frame1.data[1280] = 8'hF6; frame1.valid[1280] = 1'b1; frame1.error[1280] = 1'b0;frame1.data[1281] = 8'hF7; frame1.valid[1281] = 1'b1; frame1.error[1281] = 1'b0;frame1.data[1282] = 8'hF8; frame1.valid[1282] = 1'b1; frame1.error[1282] = 1'b0;frame1.data[1283] = 8'hF9; frame1.valid[1283] = 1'b1; frame1.error[1283] = 1'b0;frame1.data[1284] = 8'hFA; frame1.valid[1284] = 1'b1; frame1.error[1284] = 1'b0;frame1.data[1285] = 8'hFB; frame1.valid[1285] = 1'b1; frame1.error[1285] = 1'b0;frame1.data[1286] = 8'hFC; frame1.valid[1286] = 1'b1; frame1.error[1286] = 1'b0;frame1.data[1287] = 8'hFD; frame1.valid[1287] = 1'b1; frame1.error[1287] = 1'b0;frame1.data[1288] = 8'hFE; frame1.valid[1288] = 1'b1; frame1.error[1288] = 1'b0;frame1.data[1289] = 8'h00; frame1.valid[1289] = 1'b1; frame1.error[1289] = 1'b0;frame1.data[1290] = 8'h01; frame1.valid[1290] = 1'b1; frame1.error[1290] = 1'b0;frame1.data[1291] = 8'h02; frame1.valid[1291] = 1'b1; frame1.error[1291] = 1'b0;frame1.data[1292] = 8'h03; frame1.valid[1292] = 1'b1; frame1.error[1292] = 1'b0;frame1.data[1293] = 8'h04; frame1.valid[1293] = 1'b1; frame1.error[1293] = 1'b0;
        frame1.data[1294] = 8'h05; frame1.valid[1294] = 1'b1; frame1.error[1294] = 1'b0;frame1.data[1295] = 8'h06; frame1.valid[1295] = 1'b1; frame1.error[1295] = 1'b0;frame1.data[1296] = 8'h07; frame1.valid[1296] = 1'b1; frame1.error[1296] = 1'b0;frame1.data[1297] = 8'h08; frame1.valid[1297] = 1'b1; frame1.error[1297] = 1'b0;frame1.data[1298] = 8'h09; frame1.valid[1298] = 1'b1; frame1.error[1298] = 1'b0;frame1.data[1299] = 8'h0A; frame1.valid[1299] = 1'b1; frame1.error[1299] = 1'b0;frame1.data[1300] = 8'h0B; frame1.valid[1300] = 1'b1; frame1.error[1300] = 1'b0;frame1.data[1301] = 8'h0C; frame1.valid[1301] = 1'b1; frame1.error[1301] = 1'b0;frame1.data[1302] = 8'h0D; frame1.valid[1302] = 1'b1; frame1.error[1302] = 1'b0;frame1.data[1303] = 8'h0E; frame1.valid[1303] = 1'b1; frame1.error[1303] = 1'b0;frame1.data[1304] = 8'h0F; frame1.valid[1304] = 1'b1; frame1.error[1304] = 1'b0;frame1.data[1305] = 8'h10; frame1.valid[1305] = 1'b1; frame1.error[1305] = 1'b0;frame1.data[1306] = 8'h11; frame1.valid[1306] = 1'b1; frame1.error[1306] = 1'b0;frame1.data[1307] = 8'h12; frame1.valid[1307] = 1'b1; frame1.error[1307] = 1'b0;frame1.data[1308] = 8'h13; frame1.valid[1308] = 1'b1; frame1.error[1308] = 1'b0;frame1.data[1309] = 8'h14; frame1.valid[1309] = 1'b1; frame1.error[1309] = 1'b0;
        frame1.data[1310] = 8'h15; frame1.valid[1310] = 1'b1; frame1.error[1310] = 1'b0;frame1.data[1311] = 8'h16; frame1.valid[1311] = 1'b1; frame1.error[1311] = 1'b0;frame1.data[1312] = 8'h17; frame1.valid[1312] = 1'b1; frame1.error[1312] = 1'b0;frame1.data[1313] = 8'h18; frame1.valid[1313] = 1'b1; frame1.error[1313] = 1'b0;frame1.data[1314] = 8'h19; frame1.valid[1314] = 1'b1; frame1.error[1314] = 1'b0;frame1.data[1315] = 8'h1A; frame1.valid[1315] = 1'b1; frame1.error[1315] = 1'b0;frame1.data[1316] = 8'h1B; frame1.valid[1316] = 1'b1; frame1.error[1316] = 1'b0;frame1.data[1317] = 8'h1C; frame1.valid[1317] = 1'b1; frame1.error[1317] = 1'b0;frame1.data[1318] = 8'h1D; frame1.valid[1318] = 1'b1; frame1.error[1318] = 1'b0;frame1.data[1319] = 8'h1E; frame1.valid[1319] = 1'b1; frame1.error[1319] = 1'b0;frame1.data[1320] = 8'h1F; frame1.valid[1320] = 1'b1; frame1.error[1320] = 1'b0;frame1.data[1321] = 8'h20; frame1.valid[1321] = 1'b1; frame1.error[1321] = 1'b0;frame1.data[1322] = 8'h21; frame1.valid[1322] = 1'b1; frame1.error[1322] = 1'b0;frame1.data[1323] = 8'h22; frame1.valid[1323] = 1'b1; frame1.error[1323] = 1'b0;frame1.data[1324] = 8'h23; frame1.valid[1324] = 1'b1; frame1.error[1324] = 1'b0;frame1.data[1325] = 8'h24; frame1.valid[1325] = 1'b1; frame1.error[1325] = 1'b0;
        frame1.data[1326] = 8'h25; frame1.valid[1326] = 1'b1; frame1.error[1326] = 1'b0;frame1.data[1327] = 8'h26; frame1.valid[1327] = 1'b1; frame1.error[1327] = 1'b0;frame1.data[1328] = 8'h27; frame1.valid[1328] = 1'b1; frame1.error[1328] = 1'b0;frame1.data[1329] = 8'h28; frame1.valid[1329] = 1'b1; frame1.error[1329] = 1'b0;frame1.data[1330] = 8'h29; frame1.valid[1330] = 1'b1; frame1.error[1330] = 1'b0;frame1.data[1331] = 8'h2A; frame1.valid[1331] = 1'b1; frame1.error[1331] = 1'b0;frame1.data[1332] = 8'h2B; frame1.valid[1332] = 1'b1; frame1.error[1332] = 1'b0;frame1.data[1333] = 8'h2C; frame1.valid[1333] = 1'b1; frame1.error[1333] = 1'b0;frame1.data[1334] = 8'h2D; frame1.valid[1334] = 1'b1; frame1.error[1334] = 1'b0;frame1.data[1335] = 8'h2E; frame1.valid[1335] = 1'b1; frame1.error[1335] = 1'b0;frame1.data[1336] = 8'h2F; frame1.valid[1336] = 1'b1; frame1.error[1336] = 1'b0;frame1.data[1337] = 8'h30; frame1.valid[1337] = 1'b1; frame1.error[1337] = 1'b0;frame1.data[1338] = 8'h31; frame1.valid[1338] = 1'b1; frame1.error[1338] = 1'b0;frame1.data[1339] = 8'h32; frame1.valid[1339] = 1'b1; frame1.error[1339] = 1'b0;frame1.data[1340] = 8'h33; frame1.valid[1340] = 1'b1; frame1.error[1340] = 1'b0;frame1.data[1341] = 8'h34; frame1.valid[1341] = 1'b1; frame1.error[1341] = 1'b0;
        frame1.data[1342] = 8'h35; frame1.valid[1342] = 1'b1; frame1.error[1342] = 1'b0;frame1.data[1343] = 8'h36; frame1.valid[1343] = 1'b1; frame1.error[1343] = 1'b0;frame1.data[1344] = 8'h37; frame1.valid[1344] = 1'b1; frame1.error[1344] = 1'b0;frame1.data[1345] = 8'h38; frame1.valid[1345] = 1'b1; frame1.error[1345] = 1'b0;frame1.data[1346] = 8'h39; frame1.valid[1346] = 1'b1; frame1.error[1346] = 1'b0;frame1.data[1347] = 8'h3A; frame1.valid[1347] = 1'b1; frame1.error[1347] = 1'b0;frame1.data[1348] = 8'h3B; frame1.valid[1348] = 1'b1; frame1.error[1348] = 1'b0;frame1.data[1349] = 8'h3C; frame1.valid[1349] = 1'b1; frame1.error[1349] = 1'b0;frame1.data[1350] = 8'h3D; frame1.valid[1350] = 1'b1; frame1.error[1350] = 1'b0;frame1.data[1351] = 8'h3E; frame1.valid[1351] = 1'b1; frame1.error[1351] = 1'b0;frame1.data[1352] = 8'h3F; frame1.valid[1352] = 1'b1; frame1.error[1352] = 1'b0;frame1.data[1353] = 8'h40; frame1.valid[1353] = 1'b1; frame1.error[1353] = 1'b0;frame1.data[1354] = 8'h41; frame1.valid[1354] = 1'b1; frame1.error[1354] = 1'b0;frame1.data[1355] = 8'h42; frame1.valid[1355] = 1'b1; frame1.error[1355] = 1'b0;frame1.data[1356] = 8'h43; frame1.valid[1356] = 1'b1; frame1.error[1356] = 1'b0;frame1.data[1357] = 8'h44; frame1.valid[1357] = 1'b1; frame1.error[1357] = 1'b0;
        frame1.data[1358] = 8'h45; frame1.valid[1358] = 1'b1; frame1.error[1358] = 1'b0;frame1.data[1359] = 8'h46; frame1.valid[1359] = 1'b1; frame1.error[1359] = 1'b0;frame1.data[1360] = 8'h47; frame1.valid[1360] = 1'b1; frame1.error[1360] = 1'b0;frame1.data[1361] = 8'h48; frame1.valid[1361] = 1'b1; frame1.error[1361] = 1'b0;frame1.data[1362] = 8'h49; frame1.valid[1362] = 1'b1; frame1.error[1362] = 1'b0;frame1.data[1363] = 8'h4A; frame1.valid[1363] = 1'b1; frame1.error[1363] = 1'b0;frame1.data[1364] = 8'h4B; frame1.valid[1364] = 1'b1; frame1.error[1364] = 1'b0;frame1.data[1365] = 8'h4C; frame1.valid[1365] = 1'b1; frame1.error[1365] = 1'b0;frame1.data[1366] = 8'h4D; frame1.valid[1366] = 1'b1; frame1.error[1366] = 1'b0;frame1.data[1367] = 8'h4E; frame1.valid[1367] = 1'b1; frame1.error[1367] = 1'b0;frame1.data[1368] = 8'h4F; frame1.valid[1368] = 1'b1; frame1.error[1368] = 1'b0;frame1.data[1369] = 8'h50; frame1.valid[1369] = 1'b1; frame1.error[1369] = 1'b0;frame1.data[1370] = 8'h51; frame1.valid[1370] = 1'b1; frame1.error[1370] = 1'b0;frame1.data[1371] = 8'h52; frame1.valid[1371] = 1'b1; frame1.error[1371] = 1'b0;frame1.data[1372] = 8'h53; frame1.valid[1372] = 1'b1; frame1.error[1372] = 1'b0;frame1.data[1373] = 8'h54; frame1.valid[1373] = 1'b1; frame1.error[1373] = 1'b0;
        frame1.data[1374] = 8'h55; frame1.valid[1374] = 1'b1; frame1.error[1374] = 1'b0;frame1.data[1375] = 8'h56; frame1.valid[1375] = 1'b1; frame1.error[1375] = 1'b0;frame1.data[1376] = 8'h57; frame1.valid[1376] = 1'b1; frame1.error[1376] = 1'b0;frame1.data[1377] = 8'h58; frame1.valid[1377] = 1'b1; frame1.error[1377] = 1'b0;frame1.data[1378] = 8'h59; frame1.valid[1378] = 1'b1; frame1.error[1378] = 1'b0;frame1.data[1379] = 8'h5A; frame1.valid[1379] = 1'b1; frame1.error[1379] = 1'b0;frame1.data[1380] = 8'h5B; frame1.valid[1380] = 1'b1; frame1.error[1380] = 1'b0;frame1.data[1381] = 8'h5C; frame1.valid[1381] = 1'b1; frame1.error[1381] = 1'b0;frame1.data[1382] = 8'h5D; frame1.valid[1382] = 1'b1; frame1.error[1382] = 1'b0;frame1.data[1383] = 8'h5E; frame1.valid[1383] = 1'b1; frame1.error[1383] = 1'b0;frame1.data[1384] = 8'h5F; frame1.valid[1384] = 1'b1; frame1.error[1384] = 1'b0;frame1.data[1385] = 8'h60; frame1.valid[1385] = 1'b1; frame1.error[1385] = 1'b0;frame1.data[1386] = 8'h61; frame1.valid[1386] = 1'b1; frame1.error[1386] = 1'b0;frame1.data[1387] = 8'h62; frame1.valid[1387] = 1'b1; frame1.error[1387] = 1'b0;frame1.data[1388] = 8'h63; frame1.valid[1388] = 1'b1; frame1.error[1388] = 1'b0;frame1.data[1389] = 8'h64; frame1.valid[1389] = 1'b1; frame1.error[1389] = 1'b0;
        frame1.data[1390] = 8'h65; frame1.valid[1390] = 1'b1; frame1.error[1390] = 1'b0;frame1.data[1391] = 8'h66; frame1.valid[1391] = 1'b1; frame1.error[1391] = 1'b0;frame1.data[1392] = 8'h67; frame1.valid[1392] = 1'b1; frame1.error[1392] = 1'b0;frame1.data[1393] = 8'h68; frame1.valid[1393] = 1'b1; frame1.error[1393] = 1'b0;frame1.data[1394] = 8'h69; frame1.valid[1394] = 1'b1; frame1.error[1394] = 1'b0;frame1.data[1395] = 8'h6A; frame1.valid[1395] = 1'b1; frame1.error[1395] = 1'b0;frame1.data[1396] = 8'h6B; frame1.valid[1396] = 1'b1; frame1.error[1396] = 1'b0;frame1.data[1397] = 8'h6C; frame1.valid[1397] = 1'b1; frame1.error[1397] = 1'b0;frame1.data[1398] = 8'h6D; frame1.valid[1398] = 1'b1; frame1.error[1398] = 1'b0;frame1.data[1399] = 8'h6E; frame1.valid[1399] = 1'b1; frame1.error[1399] = 1'b0;frame1.data[1400] = 8'h6F; frame1.valid[1400] = 1'b1; frame1.error[1400] = 1'b0;frame1.data[1401] = 8'h70; frame1.valid[1401] = 1'b1; frame1.error[1401] = 1'b0;frame1.data[1402] = 8'h71; frame1.valid[1402] = 1'b1; frame1.error[1402] = 1'b0;frame1.data[1403] = 8'h72; frame1.valid[1403] = 1'b1; frame1.error[1403] = 1'b0;frame1.data[1404] = 8'h73; frame1.valid[1404] = 1'b1; frame1.error[1404] = 1'b0;frame1.data[1405] = 8'h74; frame1.valid[1405] = 1'b1; frame1.error[1405] = 1'b0;
        frame1.data[1406] = 8'h75; frame1.valid[1406] = 1'b1; frame1.error[1406] = 1'b0;frame1.data[1407] = 8'h76; frame1.valid[1407] = 1'b1; frame1.error[1407] = 1'b0;frame1.data[1408] = 8'h77; frame1.valid[1408] = 1'b1; frame1.error[1408] = 1'b0;frame1.data[1409] = 8'h78; frame1.valid[1409] = 1'b1; frame1.error[1409] = 1'b0;frame1.data[1410] = 8'h79; frame1.valid[1410] = 1'b1; frame1.error[1410] = 1'b0;frame1.data[1411] = 8'h7A; frame1.valid[1411] = 1'b1; frame1.error[1411] = 1'b0;frame1.data[1412] = 8'h7B; frame1.valid[1412] = 1'b1; frame1.error[1412] = 1'b0;frame1.data[1413] = 8'h7C; frame1.valid[1413] = 1'b1; frame1.error[1413] = 1'b0;frame1.data[1414] = 8'h7D; frame1.valid[1414] = 1'b1; frame1.error[1414] = 1'b0;frame1.data[1415] = 8'h7E; frame1.valid[1415] = 1'b1; frame1.error[1415] = 1'b0;frame1.data[1416] = 8'h7F; frame1.valid[1416] = 1'b1; frame1.error[1416] = 1'b0;frame1.data[1417] = 8'h80; frame1.valid[1417] = 1'b1; frame1.error[1417] = 1'b0;frame1.data[1418] = 8'h81; frame1.valid[1418] = 1'b1; frame1.error[1418] = 1'b0;frame1.data[1419] = 8'h82; frame1.valid[1419] = 1'b1; frame1.error[1419] = 1'b0;frame1.data[1420] = 8'h83; frame1.valid[1420] = 1'b1; frame1.error[1420] = 1'b0;frame1.data[1421] = 8'h84; frame1.valid[1421] = 1'b1; frame1.error[1421] = 1'b0;
        frame1.data[1422] = 8'h85; frame1.valid[1422] = 1'b1; frame1.error[1422] = 1'b0;frame1.data[1423] = 8'h86; frame1.valid[1423] = 1'b1; frame1.error[1423] = 1'b0;frame1.data[1424] = 8'h87; frame1.valid[1424] = 1'b1; frame1.error[1424] = 1'b0;frame1.data[1425] = 8'h88; frame1.valid[1425] = 1'b1; frame1.error[1425] = 1'b0;frame1.data[1426] = 8'h89; frame1.valid[1426] = 1'b1; frame1.error[1426] = 1'b0;frame1.data[1427] = 8'h8A; frame1.valid[1427] = 1'b1; frame1.error[1427] = 1'b0;frame1.data[1428] = 8'h8B; frame1.valid[1428] = 1'b1; frame1.error[1428] = 1'b0;frame1.data[1429] = 8'h8C; frame1.valid[1429] = 1'b1; frame1.error[1429] = 1'b0;frame1.data[1430] = 8'h8D; frame1.valid[1430] = 1'b1; frame1.error[1430] = 1'b0;frame1.data[1431] = 8'h8E; frame1.valid[1431] = 1'b1; frame1.error[1431] = 1'b0;frame1.data[1432] = 8'h8F; frame1.valid[1432] = 1'b1; frame1.error[1432] = 1'b0;frame1.data[1433] = 8'h90; frame1.valid[1433] = 1'b1; frame1.error[1433] = 1'b0;frame1.data[1434] = 8'h91; frame1.valid[1434] = 1'b1; frame1.error[1434] = 1'b0;frame1.data[1435] = 8'h92; frame1.valid[1435] = 1'b1; frame1.error[1435] = 1'b0;frame1.data[1436] = 8'h93; frame1.valid[1436] = 1'b1; frame1.error[1436] = 1'b0;frame1.data[1437] = 8'h94; frame1.valid[1437] = 1'b1; frame1.error[1437] = 1'b0;
        frame1.data[1438] = 8'h95; frame1.valid[1438] = 1'b1; frame1.error[1438] = 1'b0;frame1.data[1439] = 8'h96; frame1.valid[1439] = 1'b1; frame1.error[1439] = 1'b0;frame1.data[1440] = 8'h97; frame1.valid[1440] = 1'b1; frame1.error[1440] = 1'b0;frame1.data[1441] = 8'h98; frame1.valid[1441] = 1'b1; frame1.error[1441] = 1'b0;frame1.data[1442] = 8'h99; frame1.valid[1442] = 1'b1; frame1.error[1442] = 1'b0;frame1.data[1443] = 8'h9A; frame1.valid[1443] = 1'b1; frame1.error[1443] = 1'b0;frame1.data[1444] = 8'h9B; frame1.valid[1444] = 1'b1; frame1.error[1444] = 1'b0;frame1.data[1445] = 8'h9C; frame1.valid[1445] = 1'b1; frame1.error[1445] = 1'b0;frame1.data[1446] = 8'h9D; frame1.valid[1446] = 1'b1; frame1.error[1446] = 1'b0;frame1.data[1447] = 8'h9E; frame1.valid[1447] = 1'b1; frame1.error[1447] = 1'b0;frame1.data[1448] = 8'h9F; frame1.valid[1448] = 1'b1; frame1.error[1448] = 1'b0;frame1.data[1449] = 8'hA0; frame1.valid[1449] = 1'b1; frame1.error[1449] = 1'b0;frame1.data[1450] = 8'hA1; frame1.valid[1450] = 1'b1; frame1.error[1450] = 1'b0;frame1.data[1451] = 8'hA2; frame1.valid[1451] = 1'b1; frame1.error[1451] = 1'b0;frame1.data[1452] = 8'hA3; frame1.valid[1452] = 1'b1; frame1.error[1452] = 1'b0;frame1.data[1453] = 8'hA4; frame1.valid[1453] = 1'b1; frame1.error[1453] = 1'b0;
        frame1.data[1454] = 8'hA5; frame1.valid[1454] = 1'b1; frame1.error[1454] = 1'b0;frame1.data[1455] = 8'hA6; frame1.valid[1455] = 1'b1; frame1.error[1455] = 1'b0;frame1.data[1456] = 8'hA7; frame1.valid[1456] = 1'b1; frame1.error[1456] = 1'b0;frame1.data[1457] = 8'hA8; frame1.valid[1457] = 1'b1; frame1.error[1457] = 1'b0;frame1.data[1458] = 8'hA9; frame1.valid[1458] = 1'b1; frame1.error[1458] = 1'b0;frame1.data[1459] = 8'hAA; frame1.valid[1459] = 1'b1; frame1.error[1459] = 1'b0;frame1.data[1460] = 8'hAB; frame1.valid[1460] = 1'b1; frame1.error[1460] = 1'b0;frame1.data[1461] = 8'hAC; frame1.valid[1461] = 1'b1; frame1.error[1461] = 1'b0;frame1.data[1462] = 8'hAD; frame1.valid[1462] = 1'b1; frame1.error[1462] = 1'b0;frame1.data[1463] = 8'hAE; frame1.valid[1463] = 1'b1; frame1.error[1463] = 1'b0;frame1.data[1464] = 8'hAF; frame1.valid[1464] = 1'b1; frame1.error[1464] = 1'b0;frame1.data[1465] = 8'hB0; frame1.valid[1465] = 1'b1; frame1.error[1465] = 1'b0;frame1.data[1466] = 8'hB1; frame1.valid[1466] = 1'b1; frame1.error[1466] = 1'b0;frame1.data[1467] = 8'hB2; frame1.valid[1467] = 1'b1; frame1.error[1467] = 1'b0;frame1.data[1468] = 8'hB3; frame1.valid[1468] = 1'b1; frame1.error[1468] = 1'b0;frame1.data[1469] = 8'hB4; frame1.valid[1469] = 1'b1; frame1.error[1469] = 1'b0;
        frame1.data[1470] = 8'hB5; frame1.valid[1470] = 1'b1; frame1.error[1470] = 1'b0;frame1.data[1471] = 8'hB6; frame1.valid[1471] = 1'b1; frame1.error[1471] = 1'b0;frame1.data[1472] = 8'hB7; frame1.valid[1472] = 1'b1; frame1.error[1472] = 1'b0;frame1.data[1473] = 8'hB8; frame1.valid[1473] = 1'b1; frame1.error[1473] = 1'b0;frame1.data[1474] = 8'hB9; frame1.valid[1474] = 1'b1; frame1.error[1474] = 1'b0;frame1.data[1475] = 8'hBA; frame1.valid[1475] = 1'b1; frame1.error[1475] = 1'b0;frame1.data[1476] = 8'hBB; frame1.valid[1476] = 1'b1; frame1.error[1476] = 1'b0;frame1.data[1477] = 8'hBC; frame1.valid[1477] = 1'b1; frame1.error[1477] = 1'b0;frame1.data[1478] = 8'hBD; frame1.valid[1478] = 1'b1; frame1.error[1478] = 1'b0;frame1.data[1479] = 8'hBE; frame1.valid[1479] = 1'b1; frame1.error[1479] = 1'b0;frame1.data[1480] = 8'hBF; frame1.valid[1480] = 1'b1; frame1.error[1480] = 1'b0;frame1.data[1481] = 8'hC0; frame1.valid[1481] = 1'b1; frame1.error[1481] = 1'b0;frame1.data[1482] = 8'hC1; frame1.valid[1482] = 1'b1; frame1.error[1482] = 1'b0;frame1.data[1483] = 8'hC2; frame1.valid[1483] = 1'b1; frame1.error[1483] = 1'b0;frame1.data[1484] = 8'hC3; frame1.valid[1484] = 1'b1; frame1.error[1484] = 1'b0;frame1.data[1485] = 8'hC4; frame1.valid[1485] = 1'b1; frame1.error[1485] = 1'b0;
        frame1.data[1486] = 8'hC5; frame1.valid[1486] = 1'b1; frame1.error[1486] = 1'b0;frame1.data[1487] = 8'hC6; frame1.valid[1487] = 1'b1; frame1.error[1487] = 1'b0;frame1.data[1488] = 8'hC7; frame1.valid[1488] = 1'b1; frame1.error[1488] = 1'b0;frame1.data[1489] = 8'hC8; frame1.valid[1489] = 1'b1; frame1.error[1489] = 1'b0;frame1.data[1490] = 8'hC9; frame1.valid[1490] = 1'b1; frame1.error[1490] = 1'b0;frame1.data[1491] = 8'hCA; frame1.valid[1491] = 1'b1; frame1.error[1491] = 1'b0;frame1.data[1492] = 8'hCB; frame1.valid[1492] = 1'b1; frame1.error[1492] = 1'b0;frame1.data[1493] = 8'hCC; frame1.valid[1493] = 1'b1; frame1.error[1493] = 1'b0;frame1.data[1494] = 8'hCD; frame1.valid[1494] = 1'b1; frame1.error[1494] = 1'b0;frame1.data[1495] = 8'hCE; frame1.valid[1495] = 1'b1; frame1.error[1495] = 1'b0;frame1.data[1496] = 8'hCF; frame1.valid[1496] = 1'b1; frame1.error[1496] = 1'b0;frame1.data[1497] = 8'hD0; frame1.valid[1497] = 1'b1; frame1.error[1497] = 1'b0;frame1.data[1498] = 8'hD1; frame1.valid[1498] = 1'b1; frame1.error[1498] = 1'b0;frame1.data[1499] = 8'hD2; frame1.valid[1499] = 1'b1; frame1.error[1499] = 1'b0;frame1.data[1500] = 8'hD3; frame1.valid[1500] = 1'b1; frame1.error[1500] = 1'b0;frame1.data[1501] = 8'hD4; frame1.valid[1501] = 1'b1; frame1.error[1501] = 1'b0;
        frame1.data[1502] = 8'hD5; frame1.valid[1502] = 1'b1; frame1.error[1502] = 1'b0;frame1.data[1503] = 8'hD6; frame1.valid[1503] = 1'b1; frame1.error[1503] = 1'b0;frame1.data[1504] = 8'hD7; frame1.valid[1504] = 1'b1; frame1.error[1504] = 1'b0;frame1.data[1505] = 8'hD8; frame1.valid[1505] = 1'b1; frame1.error[1505] = 1'b0;frame1.data[1506] = 8'hD9; frame1.valid[1506] = 1'b1; frame1.error[1506] = 1'b0;frame1.data[1507] = 8'hDA; frame1.valid[1507] = 1'b1; frame1.error[1507] = 1'b0;frame1.data[1508] = 8'hDB; frame1.valid[1508] = 1'b1; frame1.error[1508] = 1'b0;frame1.data[1509] = 8'hDC; frame1.valid[1509] = 1'b1; frame1.error[1509] = 1'b0;frame1.data[1510] = 8'hDD; frame1.valid[1510] = 1'b1; frame1.error[1510] = 1'b0;frame1.data[1511] = 8'hDE; frame1.valid[1511] = 1'b1; frame1.error[1511] = 1'b0;frame1.data[1512] = 8'hDF; frame1.valid[1512] = 1'b1; frame1.error[1512] = 1'b0;frame1.data[1513] = 8'hE0; frame1.valid[1513] = 1'b1; frame1.error[1513] = 1'b0;


        // unused
        frame1.data[1514] = 8'h00;  frame1.valid[1514] = 1'b0;  frame1.error[1514] = 1'b0;
        frame1.data[1515] = 8'h00;  frame1.valid[1515] = 1'b0;  frame1.error[1515] = 1'b0;

        // No error in this frame
        frame1.bad_frame  = 1'b0;

        //-----------
        // Frame 2
        //-----------
        frame2.data[0]  = 8'h00;  frame2.valid[0]  = 1'b1;  frame2.error[0]  = 1'b0; // Destination Address (02)
        frame2.data[1]  = 8'h00;  frame2.valid[1]  = 1'b1;  frame2.error[1]  = 1'b0;
        frame2.data[2]  = 8'h00;  frame2.valid[2]  = 1'b1;  frame2.error[2]  = 1'b0;
        frame2.data[3]  = 8'h00;  frame2.valid[3]  = 1'b1;  frame2.error[3]  = 1'b0;
        frame2.data[4]  = 8'h00;  frame2.valid[4]  = 1'b1;  frame2.error[4]  = 1'b0;
        frame2.data[5]  = 8'h02;  frame2.valid[5]  = 1'b1;  frame2.error[5]  = 1'b0;
        frame2.data[6]  = 8'h00;  frame2.valid[6]  = 1'b1;  frame2.error[6]  = 1'b0; // Source Address  (03)
        frame2.data[7]  = 8'h00;  frame2.valid[7]  = 1'b1;  frame2.error[7]  = 1'b0;
        frame2.data[8]  = 8'h00;  frame2.valid[8]  = 1'b1;  frame2.error[8]  = 1'b0;
        frame2.data[9]  = 8'h00;  frame2.valid[9]  = 1'b1;  frame2.error[9]  = 1'b0;
        frame2.data[10] = 8'h00;  frame2.valid[10] = 1'b1;  frame2.error[10] = 1'b0;
        frame2.data[11] = 8'h03;  frame2.valid[11] = 1'b1;  frame2.error[11] = 1'b0;
        frame2.data[12] = 8'h05;  frame2.valid[12] = 1'b1;  frame2.error[12] = 1'b0;
        frame2.data[13] = 8'hDC;  frame2.valid[13] = 1'b1;  frame2.error[13] = 1'b0; // Length/Type = Length = 1500

        frame2.data[  14] = 8'h00; frame2.valid[  14] = 1'b1; frame2.error[  14] = 1'b0;frame2.data[  15] = 8'h01; frame2.valid[  15] = 1'b1; frame2.error[  15] = 1'b0;frame2.data[  16] = 8'h02; frame2.valid[  16] = 1'b1; frame2.error[  16] = 1'b0;frame2.data[  17] = 8'h03; frame2.valid[  17] = 1'b1; frame2.error[  17] = 1'b0;frame2.data[  18] = 8'h04; frame2.valid[  18] = 1'b1; frame2.error[  18] = 1'b0;frame2.data[  19] = 8'h05; frame2.valid[  19] = 1'b1; frame2.error[  19] = 1'b0;frame2.data[  20] = 8'h06; frame2.valid[  20] = 1'b1; frame2.error[  20] = 1'b0;frame2.data[  21] = 8'h07; frame2.valid[  21] = 1'b1; frame2.error[  21] = 1'b0;frame2.data[  22] = 8'h08; frame2.valid[  22] = 1'b1; frame2.error[  22] = 1'b0;frame2.data[  23] = 8'h09; frame2.valid[  23] = 1'b1; frame2.error[  23] = 1'b0;frame2.data[  24] = 8'h0A; frame2.valid[  24] = 1'b1; frame2.error[  24] = 1'b0;frame2.data[  25] = 8'h0B; frame2.valid[  25] = 1'b1; frame2.error[  25] = 1'b0;frame2.data[  26] = 8'h0C; frame2.valid[  26] = 1'b1; frame2.error[  26] = 1'b0;frame2.data[  27] = 8'h0D; frame2.valid[  27] = 1'b1; frame2.error[  27] = 1'b0;frame2.data[  28] = 8'h0E; frame2.valid[  28] = 1'b1; frame2.error[  28] = 1'b0;frame2.data[  29] = 8'h0F; frame2.valid[  29] = 1'b1; frame2.error[  29] = 1'b0;
        frame2.data[  30] = 8'h10; frame2.valid[  30] = 1'b1; frame2.error[  30] = 1'b0;frame2.data[  31] = 8'h11; frame2.valid[  31] = 1'b1; frame2.error[  31] = 1'b0;frame2.data[  32] = 8'h12; frame2.valid[  32] = 1'b1; frame2.error[  32] = 1'b0;frame2.data[  33] = 8'h13; frame2.valid[  33] = 1'b1; frame2.error[  33] = 1'b0;frame2.data[  34] = 8'h14; frame2.valid[  34] = 1'b1; frame2.error[  34] = 1'b0;frame2.data[  35] = 8'h15; frame2.valid[  35] = 1'b1; frame2.error[  35] = 1'b0;frame2.data[  36] = 8'h16; frame2.valid[  36] = 1'b1; frame2.error[  36] = 1'b0;frame2.data[  37] = 8'h17; frame2.valid[  37] = 1'b1; frame2.error[  37] = 1'b0;frame2.data[  38] = 8'h18; frame2.valid[  38] = 1'b1; frame2.error[  38] = 1'b0;frame2.data[  39] = 8'h19; frame2.valid[  39] = 1'b1; frame2.error[  39] = 1'b0;frame2.data[  40] = 8'h1A; frame2.valid[  40] = 1'b1; frame2.error[  40] = 1'b0;frame2.data[  41] = 8'h1B; frame2.valid[  41] = 1'b1; frame2.error[  41] = 1'b0;frame2.data[  42] = 8'h1C; frame2.valid[  42] = 1'b1; frame2.error[  42] = 1'b0;frame2.data[  43] = 8'h1D; frame2.valid[  43] = 1'b1; frame2.error[  43] = 1'b0;frame2.data[  44] = 8'h1E; frame2.valid[  44] = 1'b1; frame2.error[  44] = 1'b0;frame2.data[  45] = 8'h1F; frame2.valid[  45] = 1'b1; frame2.error[  45] = 1'b0;
        frame2.data[  46] = 8'h20; frame2.valid[  46] = 1'b1; frame2.error[  46] = 1'b0;frame2.data[  47] = 8'h21; frame2.valid[  47] = 1'b1; frame2.error[  47] = 1'b0;frame2.data[  48] = 8'h22; frame2.valid[  48] = 1'b1; frame2.error[  48] = 1'b0;frame2.data[  49] = 8'h23; frame2.valid[  49] = 1'b1; frame2.error[  49] = 1'b0;frame2.data[  50] = 8'h24; frame2.valid[  50] = 1'b1; frame2.error[  50] = 1'b0;frame2.data[  51] = 8'h25; frame2.valid[  51] = 1'b1; frame2.error[  51] = 1'b0;frame2.data[  52] = 8'h26; frame2.valid[  52] = 1'b1; frame2.error[  52] = 1'b0;frame2.data[  53] = 8'h27; frame2.valid[  53] = 1'b1; frame2.error[  53] = 1'b0;frame2.data[  54] = 8'h28; frame2.valid[  54] = 1'b1; frame2.error[  54] = 1'b0;frame2.data[  55] = 8'h29; frame2.valid[  55] = 1'b1; frame2.error[  55] = 1'b0;frame2.data[  56] = 8'h2A; frame2.valid[  56] = 1'b1; frame2.error[  56] = 1'b0;frame2.data[  57] = 8'h2B; frame2.valid[  57] = 1'b1; frame2.error[  57] = 1'b0;frame2.data[  58] = 8'h2C; frame2.valid[  58] = 1'b1; frame2.error[  58] = 1'b0;frame2.data[  59] = 8'h2D; frame2.valid[  59] = 1'b1; frame2.error[  59] = 1'b0;frame2.data[  60] = 8'h2E; frame2.valid[  60] = 1'b1; frame2.error[  60] = 1'b0;frame2.data[  61] = 8'h2F; frame2.valid[  61] = 1'b1; frame2.error[  61] = 1'b0;
        frame2.data[  62] = 8'h30; frame2.valid[  62] = 1'b1; frame2.error[  62] = 1'b0;frame2.data[  63] = 8'h31; frame2.valid[  63] = 1'b1; frame2.error[  63] = 1'b0;frame2.data[  64] = 8'h32; frame2.valid[  64] = 1'b1; frame2.error[  64] = 1'b0;frame2.data[  65] = 8'h33; frame2.valid[  65] = 1'b1; frame2.error[  65] = 1'b0;frame2.data[  66] = 8'h34; frame2.valid[  66] = 1'b1; frame2.error[  66] = 1'b0;frame2.data[  67] = 8'h35; frame2.valid[  67] = 1'b1; frame2.error[  67] = 1'b0;frame2.data[  68] = 8'h36; frame2.valid[  68] = 1'b1; frame2.error[  68] = 1'b0;frame2.data[  69] = 8'h37; frame2.valid[  69] = 1'b1; frame2.error[  69] = 1'b0;frame2.data[  70] = 8'h38; frame2.valid[  70] = 1'b1; frame2.error[  70] = 1'b0;frame2.data[  71] = 8'h39; frame2.valid[  71] = 1'b1; frame2.error[  71] = 1'b0;frame2.data[  72] = 8'h3A; frame2.valid[  72] = 1'b1; frame2.error[  72] = 1'b0;frame2.data[  73] = 8'h3B; frame2.valid[  73] = 1'b1; frame2.error[  73] = 1'b0;frame2.data[  74] = 8'h3C; frame2.valid[  74] = 1'b1; frame2.error[  74] = 1'b0;frame2.data[  75] = 8'h3D; frame2.valid[  75] = 1'b1; frame2.error[  75] = 1'b0;frame2.data[  76] = 8'h3E; frame2.valid[  76] = 1'b1; frame2.error[  76] = 1'b0;frame2.data[  77] = 8'h3F; frame2.valid[  77] = 1'b1; frame2.error[  77] = 1'b0;
        frame2.data[  78] = 8'h40; frame2.valid[  78] = 1'b1; frame2.error[  78] = 1'b0;frame2.data[  79] = 8'h41; frame2.valid[  79] = 1'b1; frame2.error[  79] = 1'b0;frame2.data[  80] = 8'h42; frame2.valid[  80] = 1'b1; frame2.error[  80] = 1'b0;frame2.data[  81] = 8'h43; frame2.valid[  81] = 1'b1; frame2.error[  81] = 1'b0;frame2.data[  82] = 8'h44; frame2.valid[  82] = 1'b1; frame2.error[  82] = 1'b0;frame2.data[  83] = 8'h45; frame2.valid[  83] = 1'b1; frame2.error[  83] = 1'b0;frame2.data[  84] = 8'h46; frame2.valid[  84] = 1'b1; frame2.error[  84] = 1'b0;frame2.data[  85] = 8'h47; frame2.valid[  85] = 1'b1; frame2.error[  85] = 1'b0;frame2.data[  86] = 8'h48; frame2.valid[  86] = 1'b1; frame2.error[  86] = 1'b0;frame2.data[  87] = 8'h49; frame2.valid[  87] = 1'b1; frame2.error[  87] = 1'b0;frame2.data[  88] = 8'h4A; frame2.valid[  88] = 1'b1; frame2.error[  88] = 1'b0;frame2.data[  89] = 8'h4B; frame2.valid[  89] = 1'b1; frame2.error[  89] = 1'b0;frame2.data[  90] = 8'h4C; frame2.valid[  90] = 1'b1; frame2.error[  90] = 1'b0;frame2.data[  91] = 8'h4D; frame2.valid[  91] = 1'b1; frame2.error[  91] = 1'b0;frame2.data[  92] = 8'h4E; frame2.valid[  92] = 1'b1; frame2.error[  92] = 1'b0;frame2.data[  93] = 8'h4F; frame2.valid[  93] = 1'b1; frame2.error[  93] = 1'b0;
        frame2.data[  94] = 8'h50; frame2.valid[  94] = 1'b1; frame2.error[  94] = 1'b0;frame2.data[  95] = 8'h51; frame2.valid[  95] = 1'b1; frame2.error[  95] = 1'b0;frame2.data[  96] = 8'h52; frame2.valid[  96] = 1'b1; frame2.error[  96] = 1'b0;frame2.data[  97] = 8'h53; frame2.valid[  97] = 1'b1; frame2.error[  97] = 1'b0;frame2.data[  98] = 8'h54; frame2.valid[  98] = 1'b1; frame2.error[  98] = 1'b0;frame2.data[  99] = 8'h55; frame2.valid[  99] = 1'b1; frame2.error[  99] = 1'b0;frame2.data[ 100] = 8'h56; frame2.valid[ 100] = 1'b1; frame2.error[ 100] = 1'b0;frame2.data[ 101] = 8'h57; frame2.valid[ 101] = 1'b1; frame2.error[ 101] = 1'b0;frame2.data[ 102] = 8'h58; frame2.valid[ 102] = 1'b1; frame2.error[ 102] = 1'b0;frame2.data[ 103] = 8'h59; frame2.valid[ 103] = 1'b1; frame2.error[ 103] = 1'b0;frame2.data[ 104] = 8'h5A; frame2.valid[ 104] = 1'b1; frame2.error[ 104] = 1'b0;frame2.data[ 105] = 8'h5B; frame2.valid[ 105] = 1'b1; frame2.error[ 105] = 1'b0;frame2.data[ 106] = 8'h5C; frame2.valid[ 106] = 1'b1; frame2.error[ 106] = 1'b0;frame2.data[ 107] = 8'h5D; frame2.valid[ 107] = 1'b1; frame2.error[ 107] = 1'b0;frame2.data[ 108] = 8'h5E; frame2.valid[ 108] = 1'b1; frame2.error[ 108] = 1'b0;frame2.data[ 109] = 8'h5F; frame2.valid[ 109] = 1'b1; frame2.error[ 109] = 1'b0;
        frame2.data[ 110] = 8'h60; frame2.valid[ 110] = 1'b1; frame2.error[ 110] = 1'b0;frame2.data[ 111] = 8'h61; frame2.valid[ 111] = 1'b1; frame2.error[ 111] = 1'b0;frame2.data[ 112] = 8'h62; frame2.valid[ 112] = 1'b1; frame2.error[ 112] = 1'b0;frame2.data[ 113] = 8'h63; frame2.valid[ 113] = 1'b1; frame2.error[ 113] = 1'b0;frame2.data[ 114] = 8'h64; frame2.valid[ 114] = 1'b1; frame2.error[ 114] = 1'b0;frame2.data[ 115] = 8'h65; frame2.valid[ 115] = 1'b1; frame2.error[ 115] = 1'b0;frame2.data[ 116] = 8'h66; frame2.valid[ 116] = 1'b1; frame2.error[ 116] = 1'b0;frame2.data[ 117] = 8'h67; frame2.valid[ 117] = 1'b1; frame2.error[ 117] = 1'b0;frame2.data[ 118] = 8'h68; frame2.valid[ 118] = 1'b1; frame2.error[ 118] = 1'b0;frame2.data[ 119] = 8'h69; frame2.valid[ 119] = 1'b1; frame2.error[ 119] = 1'b0;frame2.data[ 120] = 8'h6A; frame2.valid[ 120] = 1'b1; frame2.error[ 120] = 1'b0;frame2.data[ 121] = 8'h6B; frame2.valid[ 121] = 1'b1; frame2.error[ 121] = 1'b0;frame2.data[ 122] = 8'h6C; frame2.valid[ 122] = 1'b1; frame2.error[ 122] = 1'b0;frame2.data[ 123] = 8'h6D; frame2.valid[ 123] = 1'b1; frame2.error[ 123] = 1'b0;frame2.data[ 124] = 8'h6E; frame2.valid[ 124] = 1'b1; frame2.error[ 124] = 1'b0;frame2.data[ 125] = 8'h6F; frame2.valid[ 125] = 1'b1; frame2.error[ 125] = 1'b0;
        frame2.data[ 126] = 8'h70; frame2.valid[ 126] = 1'b1; frame2.error[ 126] = 1'b0;frame2.data[ 127] = 8'h71; frame2.valid[ 127] = 1'b1; frame2.error[ 127] = 1'b0;frame2.data[ 128] = 8'h72; frame2.valid[ 128] = 1'b1; frame2.error[ 128] = 1'b0;frame2.data[ 129] = 8'h73; frame2.valid[ 129] = 1'b1; frame2.error[ 129] = 1'b0;frame2.data[ 130] = 8'h74; frame2.valid[ 130] = 1'b1; frame2.error[ 130] = 1'b0;frame2.data[ 131] = 8'h75; frame2.valid[ 131] = 1'b1; frame2.error[ 131] = 1'b0;frame2.data[ 132] = 8'h76; frame2.valid[ 132] = 1'b1; frame2.error[ 132] = 1'b0;frame2.data[ 133] = 8'h77; frame2.valid[ 133] = 1'b1; frame2.error[ 133] = 1'b0;frame2.data[ 134] = 8'h78; frame2.valid[ 134] = 1'b1; frame2.error[ 134] = 1'b0;frame2.data[ 135] = 8'h79; frame2.valid[ 135] = 1'b1; frame2.error[ 135] = 1'b0;frame2.data[ 136] = 8'h7A; frame2.valid[ 136] = 1'b1; frame2.error[ 136] = 1'b0;frame2.data[ 137] = 8'h7B; frame2.valid[ 137] = 1'b1; frame2.error[ 137] = 1'b0;frame2.data[ 138] = 8'h7C; frame2.valid[ 138] = 1'b1; frame2.error[ 138] = 1'b0;frame2.data[ 139] = 8'h7D; frame2.valid[ 139] = 1'b1; frame2.error[ 139] = 1'b0;frame2.data[ 140] = 8'h7E; frame2.valid[ 140] = 1'b1; frame2.error[ 140] = 1'b0;frame2.data[ 141] = 8'h7F; frame2.valid[ 141] = 1'b1; frame2.error[ 141] = 1'b0;
        frame2.data[ 142] = 8'h80; frame2.valid[ 142] = 1'b1; frame2.error[ 142] = 1'b0;frame2.data[ 143] = 8'h81; frame2.valid[ 143] = 1'b1; frame2.error[ 143] = 1'b0;frame2.data[ 144] = 8'h82; frame2.valid[ 144] = 1'b1; frame2.error[ 144] = 1'b0;frame2.data[ 145] = 8'h83; frame2.valid[ 145] = 1'b1; frame2.error[ 145] = 1'b0;frame2.data[ 146] = 8'h84; frame2.valid[ 146] = 1'b1; frame2.error[ 146] = 1'b0;frame2.data[ 147] = 8'h85; frame2.valid[ 147] = 1'b1; frame2.error[ 147] = 1'b0;frame2.data[ 148] = 8'h86; frame2.valid[ 148] = 1'b1; frame2.error[ 148] = 1'b0;frame2.data[ 149] = 8'h87; frame2.valid[ 149] = 1'b1; frame2.error[ 149] = 1'b0;frame2.data[ 150] = 8'h88; frame2.valid[ 150] = 1'b1; frame2.error[ 150] = 1'b0;frame2.data[ 151] = 8'h89; frame2.valid[ 151] = 1'b1; frame2.error[ 151] = 1'b0;frame2.data[ 152] = 8'h8A; frame2.valid[ 152] = 1'b1; frame2.error[ 152] = 1'b0;frame2.data[ 153] = 8'h8B; frame2.valid[ 153] = 1'b1; frame2.error[ 153] = 1'b0;frame2.data[ 154] = 8'h8C; frame2.valid[ 154] = 1'b1; frame2.error[ 154] = 1'b0;frame2.data[ 155] = 8'h8D; frame2.valid[ 155] = 1'b1; frame2.error[ 155] = 1'b0;frame2.data[ 156] = 8'h8E; frame2.valid[ 156] = 1'b1; frame2.error[ 156] = 1'b0;frame2.data[ 157] = 8'h8F; frame2.valid[ 157] = 1'b1; frame2.error[ 157] = 1'b0;
        frame2.data[ 158] = 8'h90; frame2.valid[ 158] = 1'b1; frame2.error[ 158] = 1'b0;frame2.data[ 159] = 8'h91; frame2.valid[ 159] = 1'b1; frame2.error[ 159] = 1'b0;frame2.data[ 160] = 8'h92; frame2.valid[ 160] = 1'b1; frame2.error[ 160] = 1'b0;frame2.data[ 161] = 8'h93; frame2.valid[ 161] = 1'b1; frame2.error[ 161] = 1'b0;frame2.data[ 162] = 8'h94; frame2.valid[ 162] = 1'b1; frame2.error[ 162] = 1'b0;frame2.data[ 163] = 8'h95; frame2.valid[ 163] = 1'b1; frame2.error[ 163] = 1'b0;frame2.data[ 164] = 8'h96; frame2.valid[ 164] = 1'b1; frame2.error[ 164] = 1'b0;frame2.data[ 165] = 8'h97; frame2.valid[ 165] = 1'b1; frame2.error[ 165] = 1'b0;frame2.data[ 166] = 8'h98; frame2.valid[ 166] = 1'b1; frame2.error[ 166] = 1'b0;frame2.data[ 167] = 8'h99; frame2.valid[ 167] = 1'b1; frame2.error[ 167] = 1'b0;frame2.data[ 168] = 8'h9A; frame2.valid[ 168] = 1'b1; frame2.error[ 168] = 1'b0;frame2.data[ 169] = 8'h9B; frame2.valid[ 169] = 1'b1; frame2.error[ 169] = 1'b0;frame2.data[ 170] = 8'h9C; frame2.valid[ 170] = 1'b1; frame2.error[ 170] = 1'b0;frame2.data[ 171] = 8'h9D; frame2.valid[ 171] = 1'b1; frame2.error[ 171] = 1'b0;frame2.data[ 172] = 8'h9E; frame2.valid[ 172] = 1'b1; frame2.error[ 172] = 1'b0;frame2.data[ 173] = 8'h9F; frame2.valid[ 173] = 1'b1; frame2.error[ 173] = 1'b0;
        frame2.data[ 174] = 8'hA0; frame2.valid[ 174] = 1'b1; frame2.error[ 174] = 1'b0;frame2.data[ 175] = 8'hA1; frame2.valid[ 175] = 1'b1; frame2.error[ 175] = 1'b0;frame2.data[ 176] = 8'hA2; frame2.valid[ 176] = 1'b1; frame2.error[ 176] = 1'b0;frame2.data[ 177] = 8'hA3; frame2.valid[ 177] = 1'b1; frame2.error[ 177] = 1'b0;frame2.data[ 178] = 8'hA4; frame2.valid[ 178] = 1'b1; frame2.error[ 178] = 1'b0;frame2.data[ 179] = 8'hA5; frame2.valid[ 179] = 1'b1; frame2.error[ 179] = 1'b0;frame2.data[ 180] = 8'hA6; frame2.valid[ 180] = 1'b1; frame2.error[ 180] = 1'b0;frame2.data[ 181] = 8'hA7; frame2.valid[ 181] = 1'b1; frame2.error[ 181] = 1'b0;frame2.data[ 182] = 8'hA8; frame2.valid[ 182] = 1'b1; frame2.error[ 182] = 1'b0;frame2.data[ 183] = 8'hA9; frame2.valid[ 183] = 1'b1; frame2.error[ 183] = 1'b0;frame2.data[ 184] = 8'hAA; frame2.valid[ 184] = 1'b1; frame2.error[ 184] = 1'b0;frame2.data[ 185] = 8'hAB; frame2.valid[ 185] = 1'b1; frame2.error[ 185] = 1'b0;frame2.data[ 186] = 8'hAC; frame2.valid[ 186] = 1'b1; frame2.error[ 186] = 1'b0;frame2.data[ 187] = 8'hAD; frame2.valid[ 187] = 1'b1; frame2.error[ 187] = 1'b0;frame2.data[ 188] = 8'hAE; frame2.valid[ 188] = 1'b1; frame2.error[ 188] = 1'b0;frame2.data[ 189] = 8'hAF; frame2.valid[ 189] = 1'b1; frame2.error[ 189] = 1'b0;
        frame2.data[ 190] = 8'hB0; frame2.valid[ 190] = 1'b1; frame2.error[ 190] = 1'b0;frame2.data[ 191] = 8'hB1; frame2.valid[ 191] = 1'b1; frame2.error[ 191] = 1'b0;frame2.data[ 192] = 8'hB2; frame2.valid[ 192] = 1'b1; frame2.error[ 192] = 1'b0;frame2.data[ 193] = 8'hB3; frame2.valid[ 193] = 1'b1; frame2.error[ 193] = 1'b0;frame2.data[ 194] = 8'hB4; frame2.valid[ 194] = 1'b1; frame2.error[ 194] = 1'b0;frame2.data[ 195] = 8'hB5; frame2.valid[ 195] = 1'b1; frame2.error[ 195] = 1'b0;frame2.data[ 196] = 8'hB6; frame2.valid[ 196] = 1'b1; frame2.error[ 196] = 1'b0;frame2.data[ 197] = 8'hB7; frame2.valid[ 197] = 1'b1; frame2.error[ 197] = 1'b0;frame2.data[ 198] = 8'hB8; frame2.valid[ 198] = 1'b1; frame2.error[ 198] = 1'b0;frame2.data[ 199] = 8'hB9; frame2.valid[ 199] = 1'b1; frame2.error[ 199] = 1'b0;frame2.data[ 200] = 8'hBA; frame2.valid[ 200] = 1'b1; frame2.error[ 200] = 1'b0;frame2.data[ 201] = 8'hBB; frame2.valid[ 201] = 1'b1; frame2.error[ 201] = 1'b0;frame2.data[ 202] = 8'hBC; frame2.valid[ 202] = 1'b1; frame2.error[ 202] = 1'b0;frame2.data[ 203] = 8'hBD; frame2.valid[ 203] = 1'b1; frame2.error[ 203] = 1'b0;frame2.data[ 204] = 8'hBE; frame2.valid[ 204] = 1'b1; frame2.error[ 204] = 1'b0;frame2.data[ 205] = 8'hBF; frame2.valid[ 205] = 1'b1; frame2.error[ 205] = 1'b0;
        frame2.data[ 206] = 8'hC0; frame2.valid[ 206] = 1'b1; frame2.error[ 206] = 1'b0;frame2.data[ 207] = 8'hC1; frame2.valid[ 207] = 1'b1; frame2.error[ 207] = 1'b0;frame2.data[ 208] = 8'hC2; frame2.valid[ 208] = 1'b1; frame2.error[ 208] = 1'b0;frame2.data[ 209] = 8'hC3; frame2.valid[ 209] = 1'b1; frame2.error[ 209] = 1'b0;frame2.data[ 210] = 8'hC4; frame2.valid[ 210] = 1'b1; frame2.error[ 210] = 1'b0;frame2.data[ 211] = 8'hC5; frame2.valid[ 211] = 1'b1; frame2.error[ 211] = 1'b0;frame2.data[ 212] = 8'hC6; frame2.valid[ 212] = 1'b1; frame2.error[ 212] = 1'b0;frame2.data[ 213] = 8'hC7; frame2.valid[ 213] = 1'b1; frame2.error[ 213] = 1'b0;frame2.data[ 214] = 8'hC8; frame2.valid[ 214] = 1'b1; frame2.error[ 214] = 1'b0;frame2.data[ 215] = 8'hC9; frame2.valid[ 215] = 1'b1; frame2.error[ 215] = 1'b0;frame2.data[ 216] = 8'hCA; frame2.valid[ 216] = 1'b1; frame2.error[ 216] = 1'b0;frame2.data[ 217] = 8'hCB; frame2.valid[ 217] = 1'b1; frame2.error[ 217] = 1'b0;frame2.data[ 218] = 8'hCC; frame2.valid[ 218] = 1'b1; frame2.error[ 218] = 1'b0;frame2.data[ 219] = 8'hCD; frame2.valid[ 219] = 1'b1; frame2.error[ 219] = 1'b0;frame2.data[ 220] = 8'hCE; frame2.valid[ 220] = 1'b1; frame2.error[ 220] = 1'b0;frame2.data[ 221] = 8'hCF; frame2.valid[ 221] = 1'b1; frame2.error[ 221] = 1'b0;
        frame2.data[ 222] = 8'hD0; frame2.valid[ 222] = 1'b1; frame2.error[ 222] = 1'b0;frame2.data[ 223] = 8'hD1; frame2.valid[ 223] = 1'b1; frame2.error[ 223] = 1'b0;frame2.data[ 224] = 8'hD2; frame2.valid[ 224] = 1'b1; frame2.error[ 224] = 1'b0;frame2.data[ 225] = 8'hD3; frame2.valid[ 225] = 1'b1; frame2.error[ 225] = 1'b0;frame2.data[ 226] = 8'hD4; frame2.valid[ 226] = 1'b1; frame2.error[ 226] = 1'b0;frame2.data[ 227] = 8'hD5; frame2.valid[ 227] = 1'b1; frame2.error[ 227] = 1'b0;frame2.data[ 228] = 8'hD6; frame2.valid[ 228] = 1'b1; frame2.error[ 228] = 1'b0;frame2.data[ 229] = 8'hD7; frame2.valid[ 229] = 1'b1; frame2.error[ 229] = 1'b0;frame2.data[ 230] = 8'hD8; frame2.valid[ 230] = 1'b1; frame2.error[ 230] = 1'b0;frame2.data[ 231] = 8'hD9; frame2.valid[ 231] = 1'b1; frame2.error[ 231] = 1'b0;frame2.data[ 232] = 8'hDA; frame2.valid[ 232] = 1'b1; frame2.error[ 232] = 1'b0;frame2.data[ 233] = 8'hDB; frame2.valid[ 233] = 1'b1; frame2.error[ 233] = 1'b0;frame2.data[ 234] = 8'hDC; frame2.valid[ 234] = 1'b1; frame2.error[ 234] = 1'b0;frame2.data[ 235] = 8'hDD; frame2.valid[ 235] = 1'b1; frame2.error[ 235] = 1'b0;frame2.data[ 236] = 8'hDE; frame2.valid[ 236] = 1'b1; frame2.error[ 236] = 1'b0;frame2.data[ 237] = 8'hDF; frame2.valid[ 237] = 1'b1; frame2.error[ 237] = 1'b0;
        frame2.data[ 238] = 8'hE0; frame2.valid[ 238] = 1'b1; frame2.error[ 238] = 1'b0;frame2.data[ 239] = 8'hE1; frame2.valid[ 239] = 1'b1; frame2.error[ 239] = 1'b0;frame2.data[ 240] = 8'hE2; frame2.valid[ 240] = 1'b1; frame2.error[ 240] = 1'b0;frame2.data[ 241] = 8'hE3; frame2.valid[ 241] = 1'b1; frame2.error[ 241] = 1'b0;frame2.data[ 242] = 8'hE4; frame2.valid[ 242] = 1'b1; frame2.error[ 242] = 1'b0;frame2.data[ 243] = 8'hE5; frame2.valid[ 243] = 1'b1; frame2.error[ 243] = 1'b0;frame2.data[ 244] = 8'hE6; frame2.valid[ 244] = 1'b1; frame2.error[ 244] = 1'b0;frame2.data[ 245] = 8'hE7; frame2.valid[ 245] = 1'b1; frame2.error[ 245] = 1'b0;frame2.data[ 246] = 8'hE8; frame2.valid[ 246] = 1'b1; frame2.error[ 246] = 1'b0;frame2.data[ 247] = 8'hE9; frame2.valid[ 247] = 1'b1; frame2.error[ 247] = 1'b0;frame2.data[ 248] = 8'hEA; frame2.valid[ 248] = 1'b1; frame2.error[ 248] = 1'b0;frame2.data[ 249] = 8'hEB; frame2.valid[ 249] = 1'b1; frame2.error[ 249] = 1'b0;frame2.data[ 250] = 8'hEC; frame2.valid[ 250] = 1'b1; frame2.error[ 250] = 1'b0;frame2.data[ 251] = 8'hED; frame2.valid[ 251] = 1'b1; frame2.error[ 251] = 1'b0;frame2.data[ 252] = 8'hEE; frame2.valid[ 252] = 1'b1; frame2.error[ 252] = 1'b0;frame2.data[ 253] = 8'hEF; frame2.valid[ 253] = 1'b1; frame2.error[ 253] = 1'b0;
        frame2.data[ 254] = 8'hF0; frame2.valid[ 254] = 1'b1; frame2.error[ 254] = 1'b0;frame2.data[ 255] = 8'hF1; frame2.valid[ 255] = 1'b1; frame2.error[ 255] = 1'b0;frame2.data[ 256] = 8'hF2; frame2.valid[ 256] = 1'b1; frame2.error[ 256] = 1'b0;frame2.data[ 257] = 8'hF3; frame2.valid[ 257] = 1'b1; frame2.error[ 257] = 1'b0;frame2.data[ 258] = 8'hF4; frame2.valid[ 258] = 1'b1; frame2.error[ 258] = 1'b0;frame2.data[ 259] = 8'hF5; frame2.valid[ 259] = 1'b1; frame2.error[ 259] = 1'b0;frame2.data[ 260] = 8'hF6; frame2.valid[ 260] = 1'b1; frame2.error[ 260] = 1'b0;frame2.data[ 261] = 8'hF7; frame2.valid[ 261] = 1'b1; frame2.error[ 261] = 1'b0;frame2.data[ 262] = 8'hF8; frame2.valid[ 262] = 1'b1; frame2.error[ 262] = 1'b0;frame2.data[ 263] = 8'hF9; frame2.valid[ 263] = 1'b1; frame2.error[ 263] = 1'b0;frame2.data[ 264] = 8'hFA; frame2.valid[ 264] = 1'b1; frame2.error[ 264] = 1'b0;frame2.data[ 265] = 8'hFB; frame2.valid[ 265] = 1'b1; frame2.error[ 265] = 1'b0;frame2.data[ 266] = 8'hFC; frame2.valid[ 266] = 1'b1; frame2.error[ 266] = 1'b0;frame2.data[ 267] = 8'hFD; frame2.valid[ 267] = 1'b1; frame2.error[ 267] = 1'b0;frame2.data[ 268] = 8'hFE; frame2.valid[ 268] = 1'b1; frame2.error[ 268] = 1'b0;frame2.data[ 269] = 8'h00; frame2.valid[ 269] = 1'b1; frame2.error[ 269] = 1'b0;
        frame2.data[ 270] = 8'h01; frame2.valid[ 270] = 1'b1; frame2.error[ 270] = 1'b0;frame2.data[ 271] = 8'h02; frame2.valid[ 271] = 1'b1; frame2.error[ 271] = 1'b0;frame2.data[ 272] = 8'h03; frame2.valid[ 272] = 1'b1; frame2.error[ 272] = 1'b0;frame2.data[ 273] = 8'h04; frame2.valid[ 273] = 1'b1; frame2.error[ 273] = 1'b0;frame2.data[ 274] = 8'h05; frame2.valid[ 274] = 1'b1; frame2.error[ 274] = 1'b0;frame2.data[ 275] = 8'h06; frame2.valid[ 275] = 1'b1; frame2.error[ 275] = 1'b0;frame2.data[ 276] = 8'h07; frame2.valid[ 276] = 1'b1; frame2.error[ 276] = 1'b0;frame2.data[ 277] = 8'h08; frame2.valid[ 277] = 1'b1; frame2.error[ 277] = 1'b0;frame2.data[ 278] = 8'h09; frame2.valid[ 278] = 1'b1; frame2.error[ 278] = 1'b0;frame2.data[ 279] = 8'h0A; frame2.valid[ 279] = 1'b1; frame2.error[ 279] = 1'b0;frame2.data[ 280] = 8'h0B; frame2.valid[ 280] = 1'b1; frame2.error[ 280] = 1'b0;frame2.data[ 281] = 8'h0C; frame2.valid[ 281] = 1'b1; frame2.error[ 281] = 1'b0;frame2.data[ 282] = 8'h0D; frame2.valid[ 282] = 1'b1; frame2.error[ 282] = 1'b0;frame2.data[ 283] = 8'h0E; frame2.valid[ 283] = 1'b1; frame2.error[ 283] = 1'b0;frame2.data[ 284] = 8'h0F; frame2.valid[ 284] = 1'b1; frame2.error[ 284] = 1'b0;frame2.data[ 285] = 8'h10; frame2.valid[ 285] = 1'b1; frame2.error[ 285] = 1'b0;
        frame2.data[ 286] = 8'h11; frame2.valid[ 286] = 1'b1; frame2.error[ 286] = 1'b0;frame2.data[ 287] = 8'h12; frame2.valid[ 287] = 1'b1; frame2.error[ 287] = 1'b0;frame2.data[ 288] = 8'h13; frame2.valid[ 288] = 1'b1; frame2.error[ 288] = 1'b0;frame2.data[ 289] = 8'h14; frame2.valid[ 289] = 1'b1; frame2.error[ 289] = 1'b0;frame2.data[ 290] = 8'h15; frame2.valid[ 290] = 1'b1; frame2.error[ 290] = 1'b0;frame2.data[ 291] = 8'h16; frame2.valid[ 291] = 1'b1; frame2.error[ 291] = 1'b0;frame2.data[ 292] = 8'h17; frame2.valid[ 292] = 1'b1; frame2.error[ 292] = 1'b0;frame2.data[ 293] = 8'h18; frame2.valid[ 293] = 1'b1; frame2.error[ 293] = 1'b0;frame2.data[ 294] = 8'h19; frame2.valid[ 294] = 1'b1; frame2.error[ 294] = 1'b0;frame2.data[ 295] = 8'h1A; frame2.valid[ 295] = 1'b1; frame2.error[ 295] = 1'b0;frame2.data[ 296] = 8'h1B; frame2.valid[ 296] = 1'b1; frame2.error[ 296] = 1'b0;frame2.data[ 297] = 8'h1C; frame2.valid[ 297] = 1'b1; frame2.error[ 297] = 1'b0;frame2.data[ 298] = 8'h1D; frame2.valid[ 298] = 1'b1; frame2.error[ 298] = 1'b0;frame2.data[ 299] = 8'h1E; frame2.valid[ 299] = 1'b1; frame2.error[ 299] = 1'b0;frame2.data[ 300] = 8'h1F; frame2.valid[ 300] = 1'b1; frame2.error[ 300] = 1'b0;frame2.data[ 301] = 8'h20; frame2.valid[ 301] = 1'b1; frame2.error[ 301] = 1'b0;
        frame2.data[ 302] = 8'h21; frame2.valid[ 302] = 1'b1; frame2.error[ 302] = 1'b0;frame2.data[ 303] = 8'h22; frame2.valid[ 303] = 1'b1; frame2.error[ 303] = 1'b0;frame2.data[ 304] = 8'h23; frame2.valid[ 304] = 1'b1; frame2.error[ 304] = 1'b0;frame2.data[ 305] = 8'h24; frame2.valid[ 305] = 1'b1; frame2.error[ 305] = 1'b0;frame2.data[ 306] = 8'h25; frame2.valid[ 306] = 1'b1; frame2.error[ 306] = 1'b0;frame2.data[ 307] = 8'h26; frame2.valid[ 307] = 1'b1; frame2.error[ 307] = 1'b0;frame2.data[ 308] = 8'h27; frame2.valid[ 308] = 1'b1; frame2.error[ 308] = 1'b0;frame2.data[ 309] = 8'h28; frame2.valid[ 309] = 1'b1; frame2.error[ 309] = 1'b0;frame2.data[ 310] = 8'h29; frame2.valid[ 310] = 1'b1; frame2.error[ 310] = 1'b0;frame2.data[ 311] = 8'h2A; frame2.valid[ 311] = 1'b1; frame2.error[ 311] = 1'b0;frame2.data[ 312] = 8'h2B; frame2.valid[ 312] = 1'b1; frame2.error[ 312] = 1'b0;frame2.data[ 313] = 8'h2C; frame2.valid[ 313] = 1'b1; frame2.error[ 313] = 1'b0;frame2.data[ 314] = 8'h2D; frame2.valid[ 314] = 1'b1; frame2.error[ 314] = 1'b0;frame2.data[ 315] = 8'h2E; frame2.valid[ 315] = 1'b1; frame2.error[ 315] = 1'b0;frame2.data[ 316] = 8'h2F; frame2.valid[ 316] = 1'b1; frame2.error[ 316] = 1'b0;frame2.data[ 317] = 8'h30; frame2.valid[ 317] = 1'b1; frame2.error[ 317] = 1'b0;
        frame2.data[ 318] = 8'h31; frame2.valid[ 318] = 1'b1; frame2.error[ 318] = 1'b0;frame2.data[ 319] = 8'h32; frame2.valid[ 319] = 1'b1; frame2.error[ 319] = 1'b0;frame2.data[ 320] = 8'h33; frame2.valid[ 320] = 1'b1; frame2.error[ 320] = 1'b0;frame2.data[ 321] = 8'h34; frame2.valid[ 321] = 1'b1; frame2.error[ 321] = 1'b0;frame2.data[ 322] = 8'h35; frame2.valid[ 322] = 1'b1; frame2.error[ 322] = 1'b0;frame2.data[ 323] = 8'h36; frame2.valid[ 323] = 1'b1; frame2.error[ 323] = 1'b0;frame2.data[ 324] = 8'h37; frame2.valid[ 324] = 1'b1; frame2.error[ 324] = 1'b0;frame2.data[ 325] = 8'h38; frame2.valid[ 325] = 1'b1; frame2.error[ 325] = 1'b0;frame2.data[ 326] = 8'h39; frame2.valid[ 326] = 1'b1; frame2.error[ 326] = 1'b0;frame2.data[ 327] = 8'h3A; frame2.valid[ 327] = 1'b1; frame2.error[ 327] = 1'b0;frame2.data[ 328] = 8'h3B; frame2.valid[ 328] = 1'b1; frame2.error[ 328] = 1'b0;frame2.data[ 329] = 8'h3C; frame2.valid[ 329] = 1'b1; frame2.error[ 329] = 1'b0;frame2.data[ 330] = 8'h3D; frame2.valid[ 330] = 1'b1; frame2.error[ 330] = 1'b0;frame2.data[ 331] = 8'h3E; frame2.valid[ 331] = 1'b1; frame2.error[ 331] = 1'b0;frame2.data[ 332] = 8'h3F; frame2.valid[ 332] = 1'b1; frame2.error[ 332] = 1'b0;frame2.data[ 333] = 8'h40; frame2.valid[ 333] = 1'b1; frame2.error[ 333] = 1'b0;
        frame2.data[ 334] = 8'h41; frame2.valid[ 334] = 1'b1; frame2.error[ 334] = 1'b0;frame2.data[ 335] = 8'h42; frame2.valid[ 335] = 1'b1; frame2.error[ 335] = 1'b0;frame2.data[ 336] = 8'h43; frame2.valid[ 336] = 1'b1; frame2.error[ 336] = 1'b0;frame2.data[ 337] = 8'h44; frame2.valid[ 337] = 1'b1; frame2.error[ 337] = 1'b0;frame2.data[ 338] = 8'h45; frame2.valid[ 338] = 1'b1; frame2.error[ 338] = 1'b0;frame2.data[ 339] = 8'h46; frame2.valid[ 339] = 1'b1; frame2.error[ 339] = 1'b0;frame2.data[ 340] = 8'h47; frame2.valid[ 340] = 1'b1; frame2.error[ 340] = 1'b0;frame2.data[ 341] = 8'h48; frame2.valid[ 341] = 1'b1; frame2.error[ 341] = 1'b0;frame2.data[ 342] = 8'h49; frame2.valid[ 342] = 1'b1; frame2.error[ 342] = 1'b0;frame2.data[ 343] = 8'h4A; frame2.valid[ 343] = 1'b1; frame2.error[ 343] = 1'b0;frame2.data[ 344] = 8'h4B; frame2.valid[ 344] = 1'b1; frame2.error[ 344] = 1'b0;frame2.data[ 345] = 8'h4C; frame2.valid[ 345] = 1'b1; frame2.error[ 345] = 1'b0;frame2.data[ 346] = 8'h4D; frame2.valid[ 346] = 1'b1; frame2.error[ 346] = 1'b0;frame2.data[ 347] = 8'h4E; frame2.valid[ 347] = 1'b1; frame2.error[ 347] = 1'b0;frame2.data[ 348] = 8'h4F; frame2.valid[ 348] = 1'b1; frame2.error[ 348] = 1'b0;frame2.data[ 349] = 8'h50; frame2.valid[ 349] = 1'b1; frame2.error[ 349] = 1'b0;
        frame2.data[ 350] = 8'h51; frame2.valid[ 350] = 1'b1; frame2.error[ 350] = 1'b0;frame2.data[ 351] = 8'h52; frame2.valid[ 351] = 1'b1; frame2.error[ 351] = 1'b0;frame2.data[ 352] = 8'h53; frame2.valid[ 352] = 1'b1; frame2.error[ 352] = 1'b0;frame2.data[ 353] = 8'h54; frame2.valid[ 353] = 1'b1; frame2.error[ 353] = 1'b0;frame2.data[ 354] = 8'h55; frame2.valid[ 354] = 1'b1; frame2.error[ 354] = 1'b0;frame2.data[ 355] = 8'h56; frame2.valid[ 355] = 1'b1; frame2.error[ 355] = 1'b0;frame2.data[ 356] = 8'h57; frame2.valid[ 356] = 1'b1; frame2.error[ 356] = 1'b0;frame2.data[ 357] = 8'h58; frame2.valid[ 357] = 1'b1; frame2.error[ 357] = 1'b0;frame2.data[ 358] = 8'h59; frame2.valid[ 358] = 1'b1; frame2.error[ 358] = 1'b0;frame2.data[ 359] = 8'h5A; frame2.valid[ 359] = 1'b1; frame2.error[ 359] = 1'b0;frame2.data[ 360] = 8'h5B; frame2.valid[ 360] = 1'b1; frame2.error[ 360] = 1'b0;frame2.data[ 361] = 8'h5C; frame2.valid[ 361] = 1'b1; frame2.error[ 361] = 1'b0;frame2.data[ 362] = 8'h5D; frame2.valid[ 362] = 1'b1; frame2.error[ 362] = 1'b0;frame2.data[ 363] = 8'h5E; frame2.valid[ 363] = 1'b1; frame2.error[ 363] = 1'b0;frame2.data[ 364] = 8'h5F; frame2.valid[ 364] = 1'b1; frame2.error[ 364] = 1'b0;frame2.data[ 365] = 8'h60; frame2.valid[ 365] = 1'b1; frame2.error[ 365] = 1'b0;
        frame2.data[ 366] = 8'h61; frame2.valid[ 366] = 1'b1; frame2.error[ 366] = 1'b0;frame2.data[ 367] = 8'h62; frame2.valid[ 367] = 1'b1; frame2.error[ 367] = 1'b0;frame2.data[ 368] = 8'h63; frame2.valid[ 368] = 1'b1; frame2.error[ 368] = 1'b0;frame2.data[ 369] = 8'h64; frame2.valid[ 369] = 1'b1; frame2.error[ 369] = 1'b0;frame2.data[ 370] = 8'h65; frame2.valid[ 370] = 1'b1; frame2.error[ 370] = 1'b0;frame2.data[ 371] = 8'h66; frame2.valid[ 371] = 1'b1; frame2.error[ 371] = 1'b0;frame2.data[ 372] = 8'h67; frame2.valid[ 372] = 1'b1; frame2.error[ 372] = 1'b0;frame2.data[ 373] = 8'h68; frame2.valid[ 373] = 1'b1; frame2.error[ 373] = 1'b0;frame2.data[ 374] = 8'h69; frame2.valid[ 374] = 1'b1; frame2.error[ 374] = 1'b0;frame2.data[ 375] = 8'h6A; frame2.valid[ 375] = 1'b1; frame2.error[ 375] = 1'b0;frame2.data[ 376] = 8'h6B; frame2.valid[ 376] = 1'b1; frame2.error[ 376] = 1'b0;frame2.data[ 377] = 8'h6C; frame2.valid[ 377] = 1'b1; frame2.error[ 377] = 1'b0;frame2.data[ 378] = 8'h6D; frame2.valid[ 378] = 1'b1; frame2.error[ 378] = 1'b0;frame2.data[ 379] = 8'h6E; frame2.valid[ 379] = 1'b1; frame2.error[ 379] = 1'b0;frame2.data[ 380] = 8'h6F; frame2.valid[ 380] = 1'b1; frame2.error[ 380] = 1'b0;frame2.data[ 381] = 8'h70; frame2.valid[ 381] = 1'b1; frame2.error[ 381] = 1'b0;
        frame2.data[ 382] = 8'h71; frame2.valid[ 382] = 1'b1; frame2.error[ 382] = 1'b0;frame2.data[ 383] = 8'h72; frame2.valid[ 383] = 1'b1; frame2.error[ 383] = 1'b0;frame2.data[ 384] = 8'h73; frame2.valid[ 384] = 1'b1; frame2.error[ 384] = 1'b0;frame2.data[ 385] = 8'h74; frame2.valid[ 385] = 1'b1; frame2.error[ 385] = 1'b0;frame2.data[ 386] = 8'h75; frame2.valid[ 386] = 1'b1; frame2.error[ 386] = 1'b0;frame2.data[ 387] = 8'h76; frame2.valid[ 387] = 1'b1; frame2.error[ 387] = 1'b0;frame2.data[ 388] = 8'h77; frame2.valid[ 388] = 1'b1; frame2.error[ 388] = 1'b0;frame2.data[ 389] = 8'h78; frame2.valid[ 389] = 1'b1; frame2.error[ 389] = 1'b0;frame2.data[ 390] = 8'h79; frame2.valid[ 390] = 1'b1; frame2.error[ 390] = 1'b0;frame2.data[ 391] = 8'h7A; frame2.valid[ 391] = 1'b1; frame2.error[ 391] = 1'b0;frame2.data[ 392] = 8'h7B; frame2.valid[ 392] = 1'b1; frame2.error[ 392] = 1'b0;frame2.data[ 393] = 8'h7C; frame2.valid[ 393] = 1'b1; frame2.error[ 393] = 1'b0;frame2.data[ 394] = 8'h7D; frame2.valid[ 394] = 1'b1; frame2.error[ 394] = 1'b0;frame2.data[ 395] = 8'h7E; frame2.valid[ 395] = 1'b1; frame2.error[ 395] = 1'b0;frame2.data[ 396] = 8'h7F; frame2.valid[ 396] = 1'b1; frame2.error[ 396] = 1'b0;frame2.data[ 397] = 8'h80; frame2.valid[ 397] = 1'b1; frame2.error[ 397] = 1'b0;
        frame2.data[ 398] = 8'h81; frame2.valid[ 398] = 1'b1; frame2.error[ 398] = 1'b0;frame2.data[ 399] = 8'h82; frame2.valid[ 399] = 1'b1; frame2.error[ 399] = 1'b0;frame2.data[ 400] = 8'h83; frame2.valid[ 400] = 1'b1; frame2.error[ 400] = 1'b0;frame2.data[ 401] = 8'h84; frame2.valid[ 401] = 1'b1; frame2.error[ 401] = 1'b0;frame2.data[ 402] = 8'h85; frame2.valid[ 402] = 1'b1; frame2.error[ 402] = 1'b0;frame2.data[ 403] = 8'h86; frame2.valid[ 403] = 1'b1; frame2.error[ 403] = 1'b0;frame2.data[ 404] = 8'h87; frame2.valid[ 404] = 1'b1; frame2.error[ 404] = 1'b0;frame2.data[ 405] = 8'h88; frame2.valid[ 405] = 1'b1; frame2.error[ 405] = 1'b0;frame2.data[ 406] = 8'h89; frame2.valid[ 406] = 1'b1; frame2.error[ 406] = 1'b0;frame2.data[ 407] = 8'h8A; frame2.valid[ 407] = 1'b1; frame2.error[ 407] = 1'b0;frame2.data[ 408] = 8'h8B; frame2.valid[ 408] = 1'b1; frame2.error[ 408] = 1'b0;frame2.data[ 409] = 8'h8C; frame2.valid[ 409] = 1'b1; frame2.error[ 409] = 1'b0;frame2.data[ 410] = 8'h8D; frame2.valid[ 410] = 1'b1; frame2.error[ 410] = 1'b0;frame2.data[ 411] = 8'h8E; frame2.valid[ 411] = 1'b1; frame2.error[ 411] = 1'b0;frame2.data[ 412] = 8'h8F; frame2.valid[ 412] = 1'b1; frame2.error[ 412] = 1'b0;frame2.data[ 413] = 8'h90; frame2.valid[ 413] = 1'b1; frame2.error[ 413] = 1'b0;
        frame2.data[ 414] = 8'h91; frame2.valid[ 414] = 1'b1; frame2.error[ 414] = 1'b0;frame2.data[ 415] = 8'h92; frame2.valid[ 415] = 1'b1; frame2.error[ 415] = 1'b0;frame2.data[ 416] = 8'h93; frame2.valid[ 416] = 1'b1; frame2.error[ 416] = 1'b0;frame2.data[ 417] = 8'h94; frame2.valid[ 417] = 1'b1; frame2.error[ 417] = 1'b0;frame2.data[ 418] = 8'h95; frame2.valid[ 418] = 1'b1; frame2.error[ 418] = 1'b0;frame2.data[ 419] = 8'h96; frame2.valid[ 419] = 1'b1; frame2.error[ 419] = 1'b0;frame2.data[ 420] = 8'h97; frame2.valid[ 420] = 1'b1; frame2.error[ 420] = 1'b0;frame2.data[ 421] = 8'h98; frame2.valid[ 421] = 1'b1; frame2.error[ 421] = 1'b0;frame2.data[ 422] = 8'h99; frame2.valid[ 422] = 1'b1; frame2.error[ 422] = 1'b0;frame2.data[ 423] = 8'h9A; frame2.valid[ 423] = 1'b1; frame2.error[ 423] = 1'b0;frame2.data[ 424] = 8'h9B; frame2.valid[ 424] = 1'b1; frame2.error[ 424] = 1'b0;frame2.data[ 425] = 8'h9C; frame2.valid[ 425] = 1'b1; frame2.error[ 425] = 1'b0;frame2.data[ 426] = 8'h9D; frame2.valid[ 426] = 1'b1; frame2.error[ 426] = 1'b0;frame2.data[ 427] = 8'h9E; frame2.valid[ 427] = 1'b1; frame2.error[ 427] = 1'b0;frame2.data[ 428] = 8'h9F; frame2.valid[ 428] = 1'b1; frame2.error[ 428] = 1'b0;frame2.data[ 429] = 8'hA0; frame2.valid[ 429] = 1'b1; frame2.error[ 429] = 1'b0;
        frame2.data[ 430] = 8'hA1; frame2.valid[ 430] = 1'b1; frame2.error[ 430] = 1'b0;frame2.data[ 431] = 8'hA2; frame2.valid[ 431] = 1'b1; frame2.error[ 431] = 1'b0;frame2.data[ 432] = 8'hA3; frame2.valid[ 432] = 1'b1; frame2.error[ 432] = 1'b0;frame2.data[ 433] = 8'hA4; frame2.valid[ 433] = 1'b1; frame2.error[ 433] = 1'b0;frame2.data[ 434] = 8'hA5; frame2.valid[ 434] = 1'b1; frame2.error[ 434] = 1'b0;frame2.data[ 435] = 8'hA6; frame2.valid[ 435] = 1'b1; frame2.error[ 435] = 1'b0;frame2.data[ 436] = 8'hA7; frame2.valid[ 436] = 1'b1; frame2.error[ 436] = 1'b0;frame2.data[ 437] = 8'hA8; frame2.valid[ 437] = 1'b1; frame2.error[ 437] = 1'b0;frame2.data[ 438] = 8'hA9; frame2.valid[ 438] = 1'b1; frame2.error[ 438] = 1'b0;frame2.data[ 439] = 8'hAA; frame2.valid[ 439] = 1'b1; frame2.error[ 439] = 1'b0;frame2.data[ 440] = 8'hAB; frame2.valid[ 440] = 1'b1; frame2.error[ 440] = 1'b0;frame2.data[ 441] = 8'hAC; frame2.valid[ 441] = 1'b1; frame2.error[ 441] = 1'b0;frame2.data[ 442] = 8'hAD; frame2.valid[ 442] = 1'b1; frame2.error[ 442] = 1'b0;frame2.data[ 443] = 8'hAE; frame2.valid[ 443] = 1'b1; frame2.error[ 443] = 1'b0;frame2.data[ 444] = 8'hAF; frame2.valid[ 444] = 1'b1; frame2.error[ 444] = 1'b0;frame2.data[ 445] = 8'hB0; frame2.valid[ 445] = 1'b1; frame2.error[ 445] = 1'b0;
        frame2.data[ 446] = 8'hB1; frame2.valid[ 446] = 1'b1; frame2.error[ 446] = 1'b0;frame2.data[ 447] = 8'hB2; frame2.valid[ 447] = 1'b1; frame2.error[ 447] = 1'b0;frame2.data[ 448] = 8'hB3; frame2.valid[ 448] = 1'b1; frame2.error[ 448] = 1'b0;frame2.data[ 449] = 8'hB4; frame2.valid[ 449] = 1'b1; frame2.error[ 449] = 1'b0;frame2.data[ 450] = 8'hB5; frame2.valid[ 450] = 1'b1; frame2.error[ 450] = 1'b0;frame2.data[ 451] = 8'hB6; frame2.valid[ 451] = 1'b1; frame2.error[ 451] = 1'b0;frame2.data[ 452] = 8'hB7; frame2.valid[ 452] = 1'b1; frame2.error[ 452] = 1'b0;frame2.data[ 453] = 8'hB8; frame2.valid[ 453] = 1'b1; frame2.error[ 453] = 1'b0;frame2.data[ 454] = 8'hB9; frame2.valid[ 454] = 1'b1; frame2.error[ 454] = 1'b0;frame2.data[ 455] = 8'hBA; frame2.valid[ 455] = 1'b1; frame2.error[ 455] = 1'b0;frame2.data[ 456] = 8'hBB; frame2.valid[ 456] = 1'b1; frame2.error[ 456] = 1'b0;frame2.data[ 457] = 8'hBC; frame2.valid[ 457] = 1'b1; frame2.error[ 457] = 1'b0;frame2.data[ 458] = 8'hBD; frame2.valid[ 458] = 1'b1; frame2.error[ 458] = 1'b0;frame2.data[ 459] = 8'hBE; frame2.valid[ 459] = 1'b1; frame2.error[ 459] = 1'b0;frame2.data[ 460] = 8'hBF; frame2.valid[ 460] = 1'b1; frame2.error[ 460] = 1'b0;frame2.data[ 461] = 8'hC0; frame2.valid[ 461] = 1'b1; frame2.error[ 461] = 1'b0;
        frame2.data[ 462] = 8'hC1; frame2.valid[ 462] = 1'b1; frame2.error[ 462] = 1'b0;frame2.data[ 463] = 8'hC2; frame2.valid[ 463] = 1'b1; frame2.error[ 463] = 1'b0;frame2.data[ 464] = 8'hC3; frame2.valid[ 464] = 1'b1; frame2.error[ 464] = 1'b0;frame2.data[ 465] = 8'hC4; frame2.valid[ 465] = 1'b1; frame2.error[ 465] = 1'b0;frame2.data[ 466] = 8'hC5; frame2.valid[ 466] = 1'b1; frame2.error[ 466] = 1'b0;frame2.data[ 467] = 8'hC6; frame2.valid[ 467] = 1'b1; frame2.error[ 467] = 1'b0;frame2.data[ 468] = 8'hC7; frame2.valid[ 468] = 1'b1; frame2.error[ 468] = 1'b0;frame2.data[ 469] = 8'hC8; frame2.valid[ 469] = 1'b1; frame2.error[ 469] = 1'b0;frame2.data[ 470] = 8'hC9; frame2.valid[ 470] = 1'b1; frame2.error[ 470] = 1'b0;frame2.data[ 471] = 8'hCA; frame2.valid[ 471] = 1'b1; frame2.error[ 471] = 1'b0;frame2.data[ 472] = 8'hCB; frame2.valid[ 472] = 1'b1; frame2.error[ 472] = 1'b0;frame2.data[ 473] = 8'hCC; frame2.valid[ 473] = 1'b1; frame2.error[ 473] = 1'b0;frame2.data[ 474] = 8'hCD; frame2.valid[ 474] = 1'b1; frame2.error[ 474] = 1'b0;frame2.data[ 475] = 8'hCE; frame2.valid[ 475] = 1'b1; frame2.error[ 475] = 1'b0;frame2.data[ 476] = 8'hCF; frame2.valid[ 476] = 1'b1; frame2.error[ 476] = 1'b0;frame2.data[ 477] = 8'hD0; frame2.valid[ 477] = 1'b1; frame2.error[ 477] = 1'b0;
        frame2.data[ 478] = 8'hD1; frame2.valid[ 478] = 1'b1; frame2.error[ 478] = 1'b0;frame2.data[ 479] = 8'hD2; frame2.valid[ 479] = 1'b1; frame2.error[ 479] = 1'b0;frame2.data[ 480] = 8'hD3; frame2.valid[ 480] = 1'b1; frame2.error[ 480] = 1'b0;frame2.data[ 481] = 8'hD4; frame2.valid[ 481] = 1'b1; frame2.error[ 481] = 1'b0;frame2.data[ 482] = 8'hD5; frame2.valid[ 482] = 1'b1; frame2.error[ 482] = 1'b0;frame2.data[ 483] = 8'hD6; frame2.valid[ 483] = 1'b1; frame2.error[ 483] = 1'b0;frame2.data[ 484] = 8'hD7; frame2.valid[ 484] = 1'b1; frame2.error[ 484] = 1'b0;frame2.data[ 485] = 8'hD8; frame2.valid[ 485] = 1'b1; frame2.error[ 485] = 1'b0;frame2.data[ 486] = 8'hD9; frame2.valid[ 486] = 1'b1; frame2.error[ 486] = 1'b0;frame2.data[ 487] = 8'hDA; frame2.valid[ 487] = 1'b1; frame2.error[ 487] = 1'b0;frame2.data[ 488] = 8'hDB; frame2.valid[ 488] = 1'b1; frame2.error[ 488] = 1'b0;frame2.data[ 489] = 8'hDC; frame2.valid[ 489] = 1'b1; frame2.error[ 489] = 1'b0;frame2.data[ 490] = 8'hDD; frame2.valid[ 490] = 1'b1; frame2.error[ 490] = 1'b0;frame2.data[ 491] = 8'hDE; frame2.valid[ 491] = 1'b1; frame2.error[ 491] = 1'b0;frame2.data[ 492] = 8'hDF; frame2.valid[ 492] = 1'b1; frame2.error[ 492] = 1'b0;frame2.data[ 493] = 8'hE0; frame2.valid[ 493] = 1'b1; frame2.error[ 493] = 1'b0;
        frame2.data[ 494] = 8'hE1; frame2.valid[ 494] = 1'b1; frame2.error[ 494] = 1'b0;frame2.data[ 495] = 8'hE2; frame2.valid[ 495] = 1'b1; frame2.error[ 495] = 1'b0;frame2.data[ 496] = 8'hE3; frame2.valid[ 496] = 1'b1; frame2.error[ 496] = 1'b0;frame2.data[ 497] = 8'hE4; frame2.valid[ 497] = 1'b1; frame2.error[ 497] = 1'b0;frame2.data[ 498] = 8'hE5; frame2.valid[ 498] = 1'b1; frame2.error[ 498] = 1'b0;frame2.data[ 499] = 8'hE6; frame2.valid[ 499] = 1'b1; frame2.error[ 499] = 1'b0;frame2.data[ 500] = 8'hE7; frame2.valid[ 500] = 1'b1; frame2.error[ 500] = 1'b0;frame2.data[ 501] = 8'hE8; frame2.valid[ 501] = 1'b1; frame2.error[ 501] = 1'b0;frame2.data[ 502] = 8'hE9; frame2.valid[ 502] = 1'b1; frame2.error[ 502] = 1'b0;frame2.data[ 503] = 8'hEA; frame2.valid[ 503] = 1'b1; frame2.error[ 503] = 1'b0;frame2.data[ 504] = 8'hEB; frame2.valid[ 504] = 1'b1; frame2.error[ 504] = 1'b0;frame2.data[ 505] = 8'hEC; frame2.valid[ 505] = 1'b1; frame2.error[ 505] = 1'b0;frame2.data[ 506] = 8'hED; frame2.valid[ 506] = 1'b1; frame2.error[ 506] = 1'b0;frame2.data[ 507] = 8'hEE; frame2.valid[ 507] = 1'b1; frame2.error[ 507] = 1'b0;frame2.data[ 508] = 8'hEF; frame2.valid[ 508] = 1'b1; frame2.error[ 508] = 1'b0;frame2.data[ 509] = 8'hF0; frame2.valid[ 509] = 1'b1; frame2.error[ 509] = 1'b0;
        frame2.data[ 510] = 8'hF1; frame2.valid[ 510] = 1'b1; frame2.error[ 510] = 1'b0;frame2.data[ 511] = 8'hF2; frame2.valid[ 511] = 1'b1; frame2.error[ 511] = 1'b0;frame2.data[ 512] = 8'hF3; frame2.valid[ 512] = 1'b1; frame2.error[ 512] = 1'b0;frame2.data[ 513] = 8'hF4; frame2.valid[ 513] = 1'b1; frame2.error[ 513] = 1'b0;frame2.data[ 514] = 8'hF5; frame2.valid[ 514] = 1'b1; frame2.error[ 514] = 1'b0;frame2.data[ 515] = 8'hF6; frame2.valid[ 515] = 1'b1; frame2.error[ 515] = 1'b0;frame2.data[ 516] = 8'hF7; frame2.valid[ 516] = 1'b1; frame2.error[ 516] = 1'b0;frame2.data[ 517] = 8'hF8; frame2.valid[ 517] = 1'b1; frame2.error[ 517] = 1'b0;frame2.data[ 518] = 8'hF9; frame2.valid[ 518] = 1'b1; frame2.error[ 518] = 1'b0;frame2.data[ 519] = 8'hFA; frame2.valid[ 519] = 1'b1; frame2.error[ 519] = 1'b0;frame2.data[ 520] = 8'hFB; frame2.valid[ 520] = 1'b1; frame2.error[ 520] = 1'b0;frame2.data[ 521] = 8'hFC; frame2.valid[ 521] = 1'b1; frame2.error[ 521] = 1'b0;frame2.data[ 522] = 8'hFD; frame2.valid[ 522] = 1'b1; frame2.error[ 522] = 1'b0;frame2.data[ 523] = 8'hFE; frame2.valid[ 523] = 1'b1; frame2.error[ 523] = 1'b0;frame2.data[ 524] = 8'h00; frame2.valid[ 524] = 1'b1; frame2.error[ 524] = 1'b0;frame2.data[ 525] = 8'h01; frame2.valid[ 525] = 1'b1; frame2.error[ 525] = 1'b0;
        frame2.data[ 526] = 8'h02; frame2.valid[ 526] = 1'b1; frame2.error[ 526] = 1'b0;frame2.data[ 527] = 8'h03; frame2.valid[ 527] = 1'b1; frame2.error[ 527] = 1'b0;frame2.data[ 528] = 8'h04; frame2.valid[ 528] = 1'b1; frame2.error[ 528] = 1'b0;frame2.data[ 529] = 8'h05; frame2.valid[ 529] = 1'b1; frame2.error[ 529] = 1'b0;frame2.data[ 530] = 8'h06; frame2.valid[ 530] = 1'b1; frame2.error[ 530] = 1'b0;frame2.data[ 531] = 8'h07; frame2.valid[ 531] = 1'b1; frame2.error[ 531] = 1'b0;frame2.data[ 532] = 8'h08; frame2.valid[ 532] = 1'b1; frame2.error[ 532] = 1'b0;frame2.data[ 533] = 8'h09; frame2.valid[ 533] = 1'b1; frame2.error[ 533] = 1'b0;frame2.data[ 534] = 8'h0A; frame2.valid[ 534] = 1'b1; frame2.error[ 534] = 1'b0;frame2.data[ 535] = 8'h0B; frame2.valid[ 535] = 1'b1; frame2.error[ 535] = 1'b0;frame2.data[ 536] = 8'h0C; frame2.valid[ 536] = 1'b1; frame2.error[ 536] = 1'b0;frame2.data[ 537] = 8'h0D; frame2.valid[ 537] = 1'b1; frame2.error[ 537] = 1'b0;frame2.data[ 538] = 8'h0E; frame2.valid[ 538] = 1'b1; frame2.error[ 538] = 1'b0;frame2.data[ 539] = 8'h0F; frame2.valid[ 539] = 1'b1; frame2.error[ 539] = 1'b0;frame2.data[ 540] = 8'h10; frame2.valid[ 540] = 1'b1; frame2.error[ 540] = 1'b0;frame2.data[ 541] = 8'h11; frame2.valid[ 541] = 1'b1; frame2.error[ 541] = 1'b0;
        frame2.data[ 542] = 8'h12; frame2.valid[ 542] = 1'b1; frame2.error[ 542] = 1'b0;frame2.data[ 543] = 8'h13; frame2.valid[ 543] = 1'b1; frame2.error[ 543] = 1'b0;frame2.data[ 544] = 8'h14; frame2.valid[ 544] = 1'b1; frame2.error[ 544] = 1'b0;frame2.data[ 545] = 8'h15; frame2.valid[ 545] = 1'b1; frame2.error[ 545] = 1'b0;frame2.data[ 546] = 8'h16; frame2.valid[ 546] = 1'b1; frame2.error[ 546] = 1'b0;frame2.data[ 547] = 8'h17; frame2.valid[ 547] = 1'b1; frame2.error[ 547] = 1'b0;frame2.data[ 548] = 8'h18; frame2.valid[ 548] = 1'b1; frame2.error[ 548] = 1'b0;frame2.data[ 549] = 8'h19; frame2.valid[ 549] = 1'b1; frame2.error[ 549] = 1'b0;frame2.data[ 550] = 8'h1A; frame2.valid[ 550] = 1'b1; frame2.error[ 550] = 1'b0;frame2.data[ 551] = 8'h1B; frame2.valid[ 551] = 1'b1; frame2.error[ 551] = 1'b0;frame2.data[ 552] = 8'h1C; frame2.valid[ 552] = 1'b1; frame2.error[ 552] = 1'b0;frame2.data[ 553] = 8'h1D; frame2.valid[ 553] = 1'b1; frame2.error[ 553] = 1'b0;frame2.data[ 554] = 8'h1E; frame2.valid[ 554] = 1'b1; frame2.error[ 554] = 1'b0;frame2.data[ 555] = 8'h1F; frame2.valid[ 555] = 1'b1; frame2.error[ 555] = 1'b0;frame2.data[ 556] = 8'h20; frame2.valid[ 556] = 1'b1; frame2.error[ 556] = 1'b0;frame2.data[ 557] = 8'h21; frame2.valid[ 557] = 1'b1; frame2.error[ 557] = 1'b0;
        frame2.data[ 558] = 8'h22; frame2.valid[ 558] = 1'b1; frame2.error[ 558] = 1'b0;frame2.data[ 559] = 8'h23; frame2.valid[ 559] = 1'b1; frame2.error[ 559] = 1'b0;frame2.data[ 560] = 8'h24; frame2.valid[ 560] = 1'b1; frame2.error[ 560] = 1'b0;frame2.data[ 561] = 8'h25; frame2.valid[ 561] = 1'b1; frame2.error[ 561] = 1'b0;frame2.data[ 562] = 8'h26; frame2.valid[ 562] = 1'b1; frame2.error[ 562] = 1'b0;frame2.data[ 563] = 8'h27; frame2.valid[ 563] = 1'b1; frame2.error[ 563] = 1'b0;frame2.data[ 564] = 8'h28; frame2.valid[ 564] = 1'b1; frame2.error[ 564] = 1'b0;frame2.data[ 565] = 8'h29; frame2.valid[ 565] = 1'b1; frame2.error[ 565] = 1'b0;frame2.data[ 566] = 8'h2A; frame2.valid[ 566] = 1'b1; frame2.error[ 566] = 1'b0;frame2.data[ 567] = 8'h2B; frame2.valid[ 567] = 1'b1; frame2.error[ 567] = 1'b0;frame2.data[ 568] = 8'h2C; frame2.valid[ 568] = 1'b1; frame2.error[ 568] = 1'b0;frame2.data[ 569] = 8'h2D; frame2.valid[ 569] = 1'b1; frame2.error[ 569] = 1'b0;frame2.data[ 570] = 8'h2E; frame2.valid[ 570] = 1'b1; frame2.error[ 570] = 1'b0;frame2.data[ 571] = 8'h2F; frame2.valid[ 571] = 1'b1; frame2.error[ 571] = 1'b0;frame2.data[ 572] = 8'h30; frame2.valid[ 572] = 1'b1; frame2.error[ 572] = 1'b0;frame2.data[ 573] = 8'h31; frame2.valid[ 573] = 1'b1; frame2.error[ 573] = 1'b0;
        frame2.data[ 574] = 8'h32; frame2.valid[ 574] = 1'b1; frame2.error[ 574] = 1'b0;frame2.data[ 575] = 8'h33; frame2.valid[ 575] = 1'b1; frame2.error[ 575] = 1'b0;frame2.data[ 576] = 8'h34; frame2.valid[ 576] = 1'b1; frame2.error[ 576] = 1'b0;frame2.data[ 577] = 8'h35; frame2.valid[ 577] = 1'b1; frame2.error[ 577] = 1'b0;frame2.data[ 578] = 8'h36; frame2.valid[ 578] = 1'b1; frame2.error[ 578] = 1'b0;frame2.data[ 579] = 8'h37; frame2.valid[ 579] = 1'b1; frame2.error[ 579] = 1'b0;frame2.data[ 580] = 8'h38; frame2.valid[ 580] = 1'b1; frame2.error[ 580] = 1'b0;frame2.data[ 581] = 8'h39; frame2.valid[ 581] = 1'b1; frame2.error[ 581] = 1'b0;frame2.data[ 582] = 8'h3A; frame2.valid[ 582] = 1'b1; frame2.error[ 582] = 1'b0;frame2.data[ 583] = 8'h3B; frame2.valid[ 583] = 1'b1; frame2.error[ 583] = 1'b0;frame2.data[ 584] = 8'h3C; frame2.valid[ 584] = 1'b1; frame2.error[ 584] = 1'b0;frame2.data[ 585] = 8'h3D; frame2.valid[ 585] = 1'b1; frame2.error[ 585] = 1'b0;frame2.data[ 586] = 8'h3E; frame2.valid[ 586] = 1'b1; frame2.error[ 586] = 1'b0;frame2.data[ 587] = 8'h3F; frame2.valid[ 587] = 1'b1; frame2.error[ 587] = 1'b0;frame2.data[ 588] = 8'h40; frame2.valid[ 588] = 1'b1; frame2.error[ 588] = 1'b0;frame2.data[ 589] = 8'h41; frame2.valid[ 589] = 1'b1; frame2.error[ 589] = 1'b0;
        frame2.data[ 590] = 8'h42; frame2.valid[ 590] = 1'b1; frame2.error[ 590] = 1'b0;frame2.data[ 591] = 8'h43; frame2.valid[ 591] = 1'b1; frame2.error[ 591] = 1'b0;frame2.data[ 592] = 8'h44; frame2.valid[ 592] = 1'b1; frame2.error[ 592] = 1'b0;frame2.data[ 593] = 8'h45; frame2.valid[ 593] = 1'b1; frame2.error[ 593] = 1'b0;frame2.data[ 594] = 8'h46; frame2.valid[ 594] = 1'b1; frame2.error[ 594] = 1'b0;frame2.data[ 595] = 8'h47; frame2.valid[ 595] = 1'b1; frame2.error[ 595] = 1'b0;frame2.data[ 596] = 8'h48; frame2.valid[ 596] = 1'b1; frame2.error[ 596] = 1'b0;frame2.data[ 597] = 8'h49; frame2.valid[ 597] = 1'b1; frame2.error[ 597] = 1'b0;frame2.data[ 598] = 8'h4A; frame2.valid[ 598] = 1'b1; frame2.error[ 598] = 1'b0;frame2.data[ 599] = 8'h4B; frame2.valid[ 599] = 1'b1; frame2.error[ 599] = 1'b0;frame2.data[ 600] = 8'h4C; frame2.valid[ 600] = 1'b1; frame2.error[ 600] = 1'b0;frame2.data[ 601] = 8'h4D; frame2.valid[ 601] = 1'b1; frame2.error[ 601] = 1'b0;frame2.data[ 602] = 8'h4E; frame2.valid[ 602] = 1'b1; frame2.error[ 602] = 1'b0;frame2.data[ 603] = 8'h4F; frame2.valid[ 603] = 1'b1; frame2.error[ 603] = 1'b0;frame2.data[ 604] = 8'h50; frame2.valid[ 604] = 1'b1; frame2.error[ 604] = 1'b0;frame2.data[ 605] = 8'h51; frame2.valid[ 605] = 1'b1; frame2.error[ 605] = 1'b0;
        frame2.data[ 606] = 8'h52; frame2.valid[ 606] = 1'b1; frame2.error[ 606] = 1'b0;frame2.data[ 607] = 8'h53; frame2.valid[ 607] = 1'b1; frame2.error[ 607] = 1'b0;frame2.data[ 608] = 8'h54; frame2.valid[ 608] = 1'b1; frame2.error[ 608] = 1'b0;frame2.data[ 609] = 8'h55; frame2.valid[ 609] = 1'b1; frame2.error[ 609] = 1'b0;frame2.data[ 610] = 8'h56; frame2.valid[ 610] = 1'b1; frame2.error[ 610] = 1'b0;frame2.data[ 611] = 8'h57; frame2.valid[ 611] = 1'b1; frame2.error[ 611] = 1'b0;frame2.data[ 612] = 8'h58; frame2.valid[ 612] = 1'b1; frame2.error[ 612] = 1'b0;frame2.data[ 613] = 8'h59; frame2.valid[ 613] = 1'b1; frame2.error[ 613] = 1'b0;frame2.data[ 614] = 8'h5A; frame2.valid[ 614] = 1'b1; frame2.error[ 614] = 1'b0;frame2.data[ 615] = 8'h5B; frame2.valid[ 615] = 1'b1; frame2.error[ 615] = 1'b0;frame2.data[ 616] = 8'h5C; frame2.valid[ 616] = 1'b1; frame2.error[ 616] = 1'b0;frame2.data[ 617] = 8'h5D; frame2.valid[ 617] = 1'b1; frame2.error[ 617] = 1'b0;frame2.data[ 618] = 8'h5E; frame2.valid[ 618] = 1'b1; frame2.error[ 618] = 1'b0;frame2.data[ 619] = 8'h5F; frame2.valid[ 619] = 1'b1; frame2.error[ 619] = 1'b0;frame2.data[ 620] = 8'h60; frame2.valid[ 620] = 1'b1; frame2.error[ 620] = 1'b0;frame2.data[ 621] = 8'h61; frame2.valid[ 621] = 1'b1; frame2.error[ 621] = 1'b0;
        frame2.data[ 622] = 8'h62; frame2.valid[ 622] = 1'b1; frame2.error[ 622] = 1'b0;frame2.data[ 623] = 8'h63; frame2.valid[ 623] = 1'b1; frame2.error[ 623] = 1'b0;frame2.data[ 624] = 8'h64; frame2.valid[ 624] = 1'b1; frame2.error[ 624] = 1'b0;frame2.data[ 625] = 8'h65; frame2.valid[ 625] = 1'b1; frame2.error[ 625] = 1'b0;frame2.data[ 626] = 8'h66; frame2.valid[ 626] = 1'b1; frame2.error[ 626] = 1'b0;frame2.data[ 627] = 8'h67; frame2.valid[ 627] = 1'b1; frame2.error[ 627] = 1'b0;frame2.data[ 628] = 8'h68; frame2.valid[ 628] = 1'b1; frame2.error[ 628] = 1'b0;frame2.data[ 629] = 8'h69; frame2.valid[ 629] = 1'b1; frame2.error[ 629] = 1'b0;frame2.data[ 630] = 8'h6A; frame2.valid[ 630] = 1'b1; frame2.error[ 630] = 1'b0;frame2.data[ 631] = 8'h6B; frame2.valid[ 631] = 1'b1; frame2.error[ 631] = 1'b0;frame2.data[ 632] = 8'h6C; frame2.valid[ 632] = 1'b1; frame2.error[ 632] = 1'b0;frame2.data[ 633] = 8'h6D; frame2.valid[ 633] = 1'b1; frame2.error[ 633] = 1'b0;frame2.data[ 634] = 8'h6E; frame2.valid[ 634] = 1'b1; frame2.error[ 634] = 1'b0;frame2.data[ 635] = 8'h6F; frame2.valid[ 635] = 1'b1; frame2.error[ 635] = 1'b0;frame2.data[ 636] = 8'h70; frame2.valid[ 636] = 1'b1; frame2.error[ 636] = 1'b0;frame2.data[ 637] = 8'h71; frame2.valid[ 637] = 1'b1; frame2.error[ 637] = 1'b0;
        frame2.data[ 638] = 8'h72; frame2.valid[ 638] = 1'b1; frame2.error[ 638] = 1'b0;frame2.data[ 639] = 8'h73; frame2.valid[ 639] = 1'b1; frame2.error[ 639] = 1'b0;frame2.data[ 640] = 8'h74; frame2.valid[ 640] = 1'b1; frame2.error[ 640] = 1'b0;frame2.data[ 641] = 8'h75; frame2.valid[ 641] = 1'b1; frame2.error[ 641] = 1'b0;frame2.data[ 642] = 8'h76; frame2.valid[ 642] = 1'b1; frame2.error[ 642] = 1'b0;frame2.data[ 643] = 8'h77; frame2.valid[ 643] = 1'b1; frame2.error[ 643] = 1'b0;frame2.data[ 644] = 8'h78; frame2.valid[ 644] = 1'b1; frame2.error[ 644] = 1'b0;frame2.data[ 645] = 8'h79; frame2.valid[ 645] = 1'b1; frame2.error[ 645] = 1'b0;frame2.data[ 646] = 8'h7A; frame2.valid[ 646] = 1'b1; frame2.error[ 646] = 1'b0;frame2.data[ 647] = 8'h7B; frame2.valid[ 647] = 1'b1; frame2.error[ 647] = 1'b0;frame2.data[ 648] = 8'h7C; frame2.valid[ 648] = 1'b1; frame2.error[ 648] = 1'b0;frame2.data[ 649] = 8'h7D; frame2.valid[ 649] = 1'b1; frame2.error[ 649] = 1'b0;frame2.data[ 650] = 8'h7E; frame2.valid[ 650] = 1'b1; frame2.error[ 650] = 1'b0;frame2.data[ 651] = 8'h7F; frame2.valid[ 651] = 1'b1; frame2.error[ 651] = 1'b0;frame2.data[ 652] = 8'h80; frame2.valid[ 652] = 1'b1; frame2.error[ 652] = 1'b0;frame2.data[ 653] = 8'h81; frame2.valid[ 653] = 1'b1; frame2.error[ 653] = 1'b0;
        frame2.data[ 654] = 8'h82; frame2.valid[ 654] = 1'b1; frame2.error[ 654] = 1'b0;frame2.data[ 655] = 8'h83; frame2.valid[ 655] = 1'b1; frame2.error[ 655] = 1'b0;frame2.data[ 656] = 8'h84; frame2.valid[ 656] = 1'b1; frame2.error[ 656] = 1'b0;frame2.data[ 657] = 8'h85; frame2.valid[ 657] = 1'b1; frame2.error[ 657] = 1'b0;frame2.data[ 658] = 8'h86; frame2.valid[ 658] = 1'b1; frame2.error[ 658] = 1'b0;frame2.data[ 659] = 8'h87; frame2.valid[ 659] = 1'b1; frame2.error[ 659] = 1'b0;frame2.data[ 660] = 8'h88; frame2.valid[ 660] = 1'b1; frame2.error[ 660] = 1'b0;frame2.data[ 661] = 8'h89; frame2.valid[ 661] = 1'b1; frame2.error[ 661] = 1'b0;frame2.data[ 662] = 8'h8A; frame2.valid[ 662] = 1'b1; frame2.error[ 662] = 1'b0;frame2.data[ 663] = 8'h8B; frame2.valid[ 663] = 1'b1; frame2.error[ 663] = 1'b0;frame2.data[ 664] = 8'h8C; frame2.valid[ 664] = 1'b1; frame2.error[ 664] = 1'b0;frame2.data[ 665] = 8'h8D; frame2.valid[ 665] = 1'b1; frame2.error[ 665] = 1'b0;frame2.data[ 666] = 8'h8E; frame2.valid[ 666] = 1'b1; frame2.error[ 666] = 1'b0;frame2.data[ 667] = 8'h8F; frame2.valid[ 667] = 1'b1; frame2.error[ 667] = 1'b0;frame2.data[ 668] = 8'h90; frame2.valid[ 668] = 1'b1; frame2.error[ 668] = 1'b0;frame2.data[ 669] = 8'h91; frame2.valid[ 669] = 1'b1; frame2.error[ 669] = 1'b0;
        frame2.data[ 670] = 8'h92; frame2.valid[ 670] = 1'b1; frame2.error[ 670] = 1'b0;frame2.data[ 671] = 8'h93; frame2.valid[ 671] = 1'b1; frame2.error[ 671] = 1'b0;frame2.data[ 672] = 8'h94; frame2.valid[ 672] = 1'b1; frame2.error[ 672] = 1'b0;frame2.data[ 673] = 8'h95; frame2.valid[ 673] = 1'b1; frame2.error[ 673] = 1'b0;frame2.data[ 674] = 8'h96; frame2.valid[ 674] = 1'b1; frame2.error[ 674] = 1'b0;frame2.data[ 675] = 8'h97; frame2.valid[ 675] = 1'b1; frame2.error[ 675] = 1'b0;frame2.data[ 676] = 8'h98; frame2.valid[ 676] = 1'b1; frame2.error[ 676] = 1'b0;frame2.data[ 677] = 8'h99; frame2.valid[ 677] = 1'b1; frame2.error[ 677] = 1'b0;frame2.data[ 678] = 8'h9A; frame2.valid[ 678] = 1'b1; frame2.error[ 678] = 1'b0;frame2.data[ 679] = 8'h9B; frame2.valid[ 679] = 1'b1; frame2.error[ 679] = 1'b0;frame2.data[ 680] = 8'h9C; frame2.valid[ 680] = 1'b1; frame2.error[ 680] = 1'b0;frame2.data[ 681] = 8'h9D; frame2.valid[ 681] = 1'b1; frame2.error[ 681] = 1'b0;frame2.data[ 682] = 8'h9E; frame2.valid[ 682] = 1'b1; frame2.error[ 682] = 1'b0;frame2.data[ 683] = 8'h9F; frame2.valid[ 683] = 1'b1; frame2.error[ 683] = 1'b0;frame2.data[ 684] = 8'hA0; frame2.valid[ 684] = 1'b1; frame2.error[ 684] = 1'b0;frame2.data[ 685] = 8'hA1; frame2.valid[ 685] = 1'b1; frame2.error[ 685] = 1'b0;
        frame2.data[ 686] = 8'hA2; frame2.valid[ 686] = 1'b1; frame2.error[ 686] = 1'b0;frame2.data[ 687] = 8'hA3; frame2.valid[ 687] = 1'b1; frame2.error[ 687] = 1'b0;frame2.data[ 688] = 8'hA4; frame2.valid[ 688] = 1'b1; frame2.error[ 688] = 1'b0;frame2.data[ 689] = 8'hA5; frame2.valid[ 689] = 1'b1; frame2.error[ 689] = 1'b0;frame2.data[ 690] = 8'hA6; frame2.valid[ 690] = 1'b1; frame2.error[ 690] = 1'b0;frame2.data[ 691] = 8'hA7; frame2.valid[ 691] = 1'b1; frame2.error[ 691] = 1'b0;frame2.data[ 692] = 8'hA8; frame2.valid[ 692] = 1'b1; frame2.error[ 692] = 1'b0;frame2.data[ 693] = 8'hA9; frame2.valid[ 693] = 1'b1; frame2.error[ 693] = 1'b0;frame2.data[ 694] = 8'hAA; frame2.valid[ 694] = 1'b1; frame2.error[ 694] = 1'b0;frame2.data[ 695] = 8'hAB; frame2.valid[ 695] = 1'b1; frame2.error[ 695] = 1'b0;frame2.data[ 696] = 8'hAC; frame2.valid[ 696] = 1'b1; frame2.error[ 696] = 1'b0;frame2.data[ 697] = 8'hAD; frame2.valid[ 697] = 1'b1; frame2.error[ 697] = 1'b0;frame2.data[ 698] = 8'hAE; frame2.valid[ 698] = 1'b1; frame2.error[ 698] = 1'b0;frame2.data[ 699] = 8'hAF; frame2.valid[ 699] = 1'b1; frame2.error[ 699] = 1'b0;frame2.data[ 700] = 8'hB0; frame2.valid[ 700] = 1'b1; frame2.error[ 700] = 1'b0;frame2.data[ 701] = 8'hB1; frame2.valid[ 701] = 1'b1; frame2.error[ 701] = 1'b0;
        frame2.data[ 702] = 8'hB2; frame2.valid[ 702] = 1'b1; frame2.error[ 702] = 1'b0;frame2.data[ 703] = 8'hB3; frame2.valid[ 703] = 1'b1; frame2.error[ 703] = 1'b0;frame2.data[ 704] = 8'hB4; frame2.valid[ 704] = 1'b1; frame2.error[ 704] = 1'b0;frame2.data[ 705] = 8'hB5; frame2.valid[ 705] = 1'b1; frame2.error[ 705] = 1'b0;frame2.data[ 706] = 8'hB6; frame2.valid[ 706] = 1'b1; frame2.error[ 706] = 1'b0;frame2.data[ 707] = 8'hB7; frame2.valid[ 707] = 1'b1; frame2.error[ 707] = 1'b0;frame2.data[ 708] = 8'hB8; frame2.valid[ 708] = 1'b1; frame2.error[ 708] = 1'b0;frame2.data[ 709] = 8'hB9; frame2.valid[ 709] = 1'b1; frame2.error[ 709] = 1'b0;frame2.data[ 710] = 8'hBA; frame2.valid[ 710] = 1'b1; frame2.error[ 710] = 1'b0;frame2.data[ 711] = 8'hBB; frame2.valid[ 711] = 1'b1; frame2.error[ 711] = 1'b0;frame2.data[ 712] = 8'hBC; frame2.valid[ 712] = 1'b1; frame2.error[ 712] = 1'b0;frame2.data[ 713] = 8'hBD; frame2.valid[ 713] = 1'b1; frame2.error[ 713] = 1'b0;frame2.data[ 714] = 8'hBE; frame2.valid[ 714] = 1'b1; frame2.error[ 714] = 1'b0;frame2.data[ 715] = 8'hBF; frame2.valid[ 715] = 1'b1; frame2.error[ 715] = 1'b0;frame2.data[ 716] = 8'hC0; frame2.valid[ 716] = 1'b1; frame2.error[ 716] = 1'b0;frame2.data[ 717] = 8'hC1; frame2.valid[ 717] = 1'b1; frame2.error[ 717] = 1'b0;
        frame2.data[ 718] = 8'hC2; frame2.valid[ 718] = 1'b1; frame2.error[ 718] = 1'b0;frame2.data[ 719] = 8'hC3; frame2.valid[ 719] = 1'b1; frame2.error[ 719] = 1'b0;frame2.data[ 720] = 8'hC4; frame2.valid[ 720] = 1'b1; frame2.error[ 720] = 1'b0;frame2.data[ 721] = 8'hC5; frame2.valid[ 721] = 1'b1; frame2.error[ 721] = 1'b0;frame2.data[ 722] = 8'hC6; frame2.valid[ 722] = 1'b1; frame2.error[ 722] = 1'b0;frame2.data[ 723] = 8'hC7; frame2.valid[ 723] = 1'b1; frame2.error[ 723] = 1'b0;frame2.data[ 724] = 8'hC8; frame2.valid[ 724] = 1'b1; frame2.error[ 724] = 1'b0;frame2.data[ 725] = 8'hC9; frame2.valid[ 725] = 1'b1; frame2.error[ 725] = 1'b0;frame2.data[ 726] = 8'hCA; frame2.valid[ 726] = 1'b1; frame2.error[ 726] = 1'b0;frame2.data[ 727] = 8'hCB; frame2.valid[ 727] = 1'b1; frame2.error[ 727] = 1'b0;frame2.data[ 728] = 8'hCC; frame2.valid[ 728] = 1'b1; frame2.error[ 728] = 1'b0;frame2.data[ 729] = 8'hCD; frame2.valid[ 729] = 1'b1; frame2.error[ 729] = 1'b0;frame2.data[ 730] = 8'hCE; frame2.valid[ 730] = 1'b1; frame2.error[ 730] = 1'b0;frame2.data[ 731] = 8'hCF; frame2.valid[ 731] = 1'b1; frame2.error[ 731] = 1'b0;frame2.data[ 732] = 8'hD0; frame2.valid[ 732] = 1'b1; frame2.error[ 732] = 1'b0;frame2.data[ 733] = 8'hD1; frame2.valid[ 733] = 1'b1; frame2.error[ 733] = 1'b0;
        frame2.data[ 734] = 8'hD2; frame2.valid[ 734] = 1'b1; frame2.error[ 734] = 1'b0;frame2.data[ 735] = 8'hD3; frame2.valid[ 735] = 1'b1; frame2.error[ 735] = 1'b0;frame2.data[ 736] = 8'hD4; frame2.valid[ 736] = 1'b1; frame2.error[ 736] = 1'b0;frame2.data[ 737] = 8'hD5; frame2.valid[ 737] = 1'b1; frame2.error[ 737] = 1'b0;frame2.data[ 738] = 8'hD6; frame2.valid[ 738] = 1'b1; frame2.error[ 738] = 1'b0;frame2.data[ 739] = 8'hD7; frame2.valid[ 739] = 1'b1; frame2.error[ 739] = 1'b0;frame2.data[ 740] = 8'hD8; frame2.valid[ 740] = 1'b1; frame2.error[ 740] = 1'b0;frame2.data[ 741] = 8'hD9; frame2.valid[ 741] = 1'b1; frame2.error[ 741] = 1'b0;frame2.data[ 742] = 8'hDA; frame2.valid[ 742] = 1'b1; frame2.error[ 742] = 1'b0;frame2.data[ 743] = 8'hDB; frame2.valid[ 743] = 1'b1; frame2.error[ 743] = 1'b0;frame2.data[ 744] = 8'hDC; frame2.valid[ 744] = 1'b1; frame2.error[ 744] = 1'b0;frame2.data[ 745] = 8'hDD; frame2.valid[ 745] = 1'b1; frame2.error[ 745] = 1'b0;frame2.data[ 746] = 8'hDE; frame2.valid[ 746] = 1'b1; frame2.error[ 746] = 1'b0;frame2.data[ 747] = 8'hDF; frame2.valid[ 747] = 1'b1; frame2.error[ 747] = 1'b0;frame2.data[ 748] = 8'hE0; frame2.valid[ 748] = 1'b1; frame2.error[ 748] = 1'b0;frame2.data[ 749] = 8'hE1; frame2.valid[ 749] = 1'b1; frame2.error[ 749] = 1'b0;
        frame2.data[ 750] = 8'hE2; frame2.valid[ 750] = 1'b1; frame2.error[ 750] = 1'b0;frame2.data[ 751] = 8'hE3; frame2.valid[ 751] = 1'b1; frame2.error[ 751] = 1'b0;frame2.data[ 752] = 8'hE4; frame2.valid[ 752] = 1'b1; frame2.error[ 752] = 1'b0;frame2.data[ 753] = 8'hE5; frame2.valid[ 753] = 1'b1; frame2.error[ 753] = 1'b0;frame2.data[ 754] = 8'hE6; frame2.valid[ 754] = 1'b1; frame2.error[ 754] = 1'b0;frame2.data[ 755] = 8'hE7; frame2.valid[ 755] = 1'b1; frame2.error[ 755] = 1'b0;frame2.data[ 756] = 8'hE8; frame2.valid[ 756] = 1'b1; frame2.error[ 756] = 1'b0;frame2.data[ 757] = 8'hE9; frame2.valid[ 757] = 1'b1; frame2.error[ 757] = 1'b0;frame2.data[ 758] = 8'hEA; frame2.valid[ 758] = 1'b1; frame2.error[ 758] = 1'b0;frame2.data[ 759] = 8'hEB; frame2.valid[ 759] = 1'b1; frame2.error[ 759] = 1'b0;frame2.data[ 760] = 8'hEC; frame2.valid[ 760] = 1'b1; frame2.error[ 760] = 1'b0;frame2.data[ 761] = 8'hED; frame2.valid[ 761] = 1'b1; frame2.error[ 761] = 1'b0;frame2.data[ 762] = 8'hEE; frame2.valid[ 762] = 1'b1; frame2.error[ 762] = 1'b0;frame2.data[ 763] = 8'hEF; frame2.valid[ 763] = 1'b1; frame2.error[ 763] = 1'b0;frame2.data[ 764] = 8'hF0; frame2.valid[ 764] = 1'b1; frame2.error[ 764] = 1'b0;frame2.data[ 765] = 8'hF1; frame2.valid[ 765] = 1'b1; frame2.error[ 765] = 1'b0;
        frame2.data[ 766] = 8'hF2; frame2.valid[ 766] = 1'b1; frame2.error[ 766] = 1'b0;frame2.data[ 767] = 8'hF3; frame2.valid[ 767] = 1'b1; frame2.error[ 767] = 1'b0;frame2.data[ 768] = 8'hF4; frame2.valid[ 768] = 1'b1; frame2.error[ 768] = 1'b0;frame2.data[ 769] = 8'hF5; frame2.valid[ 769] = 1'b1; frame2.error[ 769] = 1'b0;frame2.data[ 770] = 8'hF6; frame2.valid[ 770] = 1'b1; frame2.error[ 770] = 1'b0;frame2.data[ 771] = 8'hF7; frame2.valid[ 771] = 1'b1; frame2.error[ 771] = 1'b0;frame2.data[ 772] = 8'hF8; frame2.valid[ 772] = 1'b1; frame2.error[ 772] = 1'b0;frame2.data[ 773] = 8'hF9; frame2.valid[ 773] = 1'b1; frame2.error[ 773] = 1'b0;frame2.data[ 774] = 8'hFA; frame2.valid[ 774] = 1'b1; frame2.error[ 774] = 1'b0;frame2.data[ 775] = 8'hFB; frame2.valid[ 775] = 1'b1; frame2.error[ 775] = 1'b0;frame2.data[ 776] = 8'hFC; frame2.valid[ 776] = 1'b1; frame2.error[ 776] = 1'b0;frame2.data[ 777] = 8'hFD; frame2.valid[ 777] = 1'b1; frame2.error[ 777] = 1'b0;frame2.data[ 778] = 8'hFE; frame2.valid[ 778] = 1'b1; frame2.error[ 778] = 1'b0;frame2.data[ 779] = 8'h00; frame2.valid[ 779] = 1'b1; frame2.error[ 779] = 1'b0;frame2.data[ 780] = 8'h01; frame2.valid[ 780] = 1'b1; frame2.error[ 780] = 1'b0;frame2.data[ 781] = 8'h02; frame2.valid[ 781] = 1'b1; frame2.error[ 781] = 1'b0;
        frame2.data[ 782] = 8'h03; frame2.valid[ 782] = 1'b1; frame2.error[ 782] = 1'b0;frame2.data[ 783] = 8'h04; frame2.valid[ 783] = 1'b1; frame2.error[ 783] = 1'b0;frame2.data[ 784] = 8'h05; frame2.valid[ 784] = 1'b1; frame2.error[ 784] = 1'b0;frame2.data[ 785] = 8'h06; frame2.valid[ 785] = 1'b1; frame2.error[ 785] = 1'b0;frame2.data[ 786] = 8'h07; frame2.valid[ 786] = 1'b1; frame2.error[ 786] = 1'b0;frame2.data[ 787] = 8'h08; frame2.valid[ 787] = 1'b1; frame2.error[ 787] = 1'b0;frame2.data[ 788] = 8'h09; frame2.valid[ 788] = 1'b1; frame2.error[ 788] = 1'b0;frame2.data[ 789] = 8'h0A; frame2.valid[ 789] = 1'b1; frame2.error[ 789] = 1'b0;frame2.data[ 790] = 8'h0B; frame2.valid[ 790] = 1'b1; frame2.error[ 790] = 1'b0;frame2.data[ 791] = 8'h0C; frame2.valid[ 791] = 1'b1; frame2.error[ 791] = 1'b0;frame2.data[ 792] = 8'h0D; frame2.valid[ 792] = 1'b1; frame2.error[ 792] = 1'b0;frame2.data[ 793] = 8'h0E; frame2.valid[ 793] = 1'b1; frame2.error[ 793] = 1'b0;frame2.data[ 794] = 8'h0F; frame2.valid[ 794] = 1'b1; frame2.error[ 794] = 1'b0;frame2.data[ 795] = 8'h10; frame2.valid[ 795] = 1'b1; frame2.error[ 795] = 1'b0;frame2.data[ 796] = 8'h11; frame2.valid[ 796] = 1'b1; frame2.error[ 796] = 1'b0;frame2.data[ 797] = 8'h12; frame2.valid[ 797] = 1'b1; frame2.error[ 797] = 1'b0;
        frame2.data[ 798] = 8'h13; frame2.valid[ 798] = 1'b1; frame2.error[ 798] = 1'b0;frame2.data[ 799] = 8'h14; frame2.valid[ 799] = 1'b1; frame2.error[ 799] = 1'b0;frame2.data[ 800] = 8'h15; frame2.valid[ 800] = 1'b1; frame2.error[ 800] = 1'b0;frame2.data[ 801] = 8'h16; frame2.valid[ 801] = 1'b1; frame2.error[ 801] = 1'b0;frame2.data[ 802] = 8'h17; frame2.valid[ 802] = 1'b1; frame2.error[ 802] = 1'b0;frame2.data[ 803] = 8'h18; frame2.valid[ 803] = 1'b1; frame2.error[ 803] = 1'b0;frame2.data[ 804] = 8'h19; frame2.valid[ 804] = 1'b1; frame2.error[ 804] = 1'b0;frame2.data[ 805] = 8'h1A; frame2.valid[ 805] = 1'b1; frame2.error[ 805] = 1'b0;frame2.data[ 806] = 8'h1B; frame2.valid[ 806] = 1'b1; frame2.error[ 806] = 1'b0;frame2.data[ 807] = 8'h1C; frame2.valid[ 807] = 1'b1; frame2.error[ 807] = 1'b0;frame2.data[ 808] = 8'h1D; frame2.valid[ 808] = 1'b1; frame2.error[ 808] = 1'b0;frame2.data[ 809] = 8'h1E; frame2.valid[ 809] = 1'b1; frame2.error[ 809] = 1'b0;frame2.data[ 810] = 8'h1F; frame2.valid[ 810] = 1'b1; frame2.error[ 810] = 1'b0;frame2.data[ 811] = 8'h20; frame2.valid[ 811] = 1'b1; frame2.error[ 811] = 1'b0;frame2.data[ 812] = 8'h21; frame2.valid[ 812] = 1'b1; frame2.error[ 812] = 1'b0;frame2.data[ 813] = 8'h22; frame2.valid[ 813] = 1'b1; frame2.error[ 813] = 1'b0;
        frame2.data[ 814] = 8'h23; frame2.valid[ 814] = 1'b1; frame2.error[ 814] = 1'b0;frame2.data[ 815] = 8'h24; frame2.valid[ 815] = 1'b1; frame2.error[ 815] = 1'b0;frame2.data[ 816] = 8'h25; frame2.valid[ 816] = 1'b1; frame2.error[ 816] = 1'b0;frame2.data[ 817] = 8'h26; frame2.valid[ 817] = 1'b1; frame2.error[ 817] = 1'b0;frame2.data[ 818] = 8'h27; frame2.valid[ 818] = 1'b1; frame2.error[ 818] = 1'b0;frame2.data[ 819] = 8'h28; frame2.valid[ 819] = 1'b1; frame2.error[ 819] = 1'b0;frame2.data[ 820] = 8'h29; frame2.valid[ 820] = 1'b1; frame2.error[ 820] = 1'b0;frame2.data[ 821] = 8'h2A; frame2.valid[ 821] = 1'b1; frame2.error[ 821] = 1'b0;frame2.data[ 822] = 8'h2B; frame2.valid[ 822] = 1'b1; frame2.error[ 822] = 1'b0;frame2.data[ 823] = 8'h2C; frame2.valid[ 823] = 1'b1; frame2.error[ 823] = 1'b0;frame2.data[ 824] = 8'h2D; frame2.valid[ 824] = 1'b1; frame2.error[ 824] = 1'b0;frame2.data[ 825] = 8'h2E; frame2.valid[ 825] = 1'b1; frame2.error[ 825] = 1'b0;frame2.data[ 826] = 8'h2F; frame2.valid[ 826] = 1'b1; frame2.error[ 826] = 1'b0;frame2.data[ 827] = 8'h30; frame2.valid[ 827] = 1'b1; frame2.error[ 827] = 1'b0;frame2.data[ 828] = 8'h31; frame2.valid[ 828] = 1'b1; frame2.error[ 828] = 1'b0;frame2.data[ 829] = 8'h32; frame2.valid[ 829] = 1'b1; frame2.error[ 829] = 1'b0;
        frame2.data[ 830] = 8'h33; frame2.valid[ 830] = 1'b1; frame2.error[ 830] = 1'b0;frame2.data[ 831] = 8'h34; frame2.valid[ 831] = 1'b1; frame2.error[ 831] = 1'b0;frame2.data[ 832] = 8'h35; frame2.valid[ 832] = 1'b1; frame2.error[ 832] = 1'b0;frame2.data[ 833] = 8'h36; frame2.valid[ 833] = 1'b1; frame2.error[ 833] = 1'b0;frame2.data[ 834] = 8'h37; frame2.valid[ 834] = 1'b1; frame2.error[ 834] = 1'b0;frame2.data[ 835] = 8'h38; frame2.valid[ 835] = 1'b1; frame2.error[ 835] = 1'b0;frame2.data[ 836] = 8'h39; frame2.valid[ 836] = 1'b1; frame2.error[ 836] = 1'b0;frame2.data[ 837] = 8'h3A; frame2.valid[ 837] = 1'b1; frame2.error[ 837] = 1'b0;frame2.data[ 838] = 8'h3B; frame2.valid[ 838] = 1'b1; frame2.error[ 838] = 1'b0;frame2.data[ 839] = 8'h3C; frame2.valid[ 839] = 1'b1; frame2.error[ 839] = 1'b0;frame2.data[ 840] = 8'h3D; frame2.valid[ 840] = 1'b1; frame2.error[ 840] = 1'b0;frame2.data[ 841] = 8'h3E; frame2.valid[ 841] = 1'b1; frame2.error[ 841] = 1'b0;frame2.data[ 842] = 8'h3F; frame2.valid[ 842] = 1'b1; frame2.error[ 842] = 1'b0;frame2.data[ 843] = 8'h40; frame2.valid[ 843] = 1'b1; frame2.error[ 843] = 1'b0;frame2.data[ 844] = 8'h41; frame2.valid[ 844] = 1'b1; frame2.error[ 844] = 1'b0;frame2.data[ 845] = 8'h42; frame2.valid[ 845] = 1'b1; frame2.error[ 845] = 1'b0;
        frame2.data[ 846] = 8'h43; frame2.valid[ 846] = 1'b1; frame2.error[ 846] = 1'b0;frame2.data[ 847] = 8'h44; frame2.valid[ 847] = 1'b1; frame2.error[ 847] = 1'b0;frame2.data[ 848] = 8'h45; frame2.valid[ 848] = 1'b1; frame2.error[ 848] = 1'b0;frame2.data[ 849] = 8'h46; frame2.valid[ 849] = 1'b1; frame2.error[ 849] = 1'b0;frame2.data[ 850] = 8'h47; frame2.valid[ 850] = 1'b1; frame2.error[ 850] = 1'b0;frame2.data[ 851] = 8'h48; frame2.valid[ 851] = 1'b1; frame2.error[ 851] = 1'b0;frame2.data[ 852] = 8'h49; frame2.valid[ 852] = 1'b1; frame2.error[ 852] = 1'b0;frame2.data[ 853] = 8'h4A; frame2.valid[ 853] = 1'b1; frame2.error[ 853] = 1'b0;frame2.data[ 854] = 8'h4B; frame2.valid[ 854] = 1'b1; frame2.error[ 854] = 1'b0;frame2.data[ 855] = 8'h4C; frame2.valid[ 855] = 1'b1; frame2.error[ 855] = 1'b0;frame2.data[ 856] = 8'h4D; frame2.valid[ 856] = 1'b1; frame2.error[ 856] = 1'b0;frame2.data[ 857] = 8'h4E; frame2.valid[ 857] = 1'b1; frame2.error[ 857] = 1'b0;frame2.data[ 858] = 8'h4F; frame2.valid[ 858] = 1'b1; frame2.error[ 858] = 1'b0;frame2.data[ 859] = 8'h50; frame2.valid[ 859] = 1'b1; frame2.error[ 859] = 1'b0;frame2.data[ 860] = 8'h51; frame2.valid[ 860] = 1'b1; frame2.error[ 860] = 1'b0;frame2.data[ 861] = 8'h52; frame2.valid[ 861] = 1'b1; frame2.error[ 861] = 1'b0;
        frame2.data[ 862] = 8'h53; frame2.valid[ 862] = 1'b1; frame2.error[ 862] = 1'b0;frame2.data[ 863] = 8'h54; frame2.valid[ 863] = 1'b1; frame2.error[ 863] = 1'b0;frame2.data[ 864] = 8'h55; frame2.valid[ 864] = 1'b1; frame2.error[ 864] = 1'b0;frame2.data[ 865] = 8'h56; frame2.valid[ 865] = 1'b1; frame2.error[ 865] = 1'b0;frame2.data[ 866] = 8'h57; frame2.valid[ 866] = 1'b1; frame2.error[ 866] = 1'b0;frame2.data[ 867] = 8'h58; frame2.valid[ 867] = 1'b1; frame2.error[ 867] = 1'b0;frame2.data[ 868] = 8'h59; frame2.valid[ 868] = 1'b1; frame2.error[ 868] = 1'b0;frame2.data[ 869] = 8'h5A; frame2.valid[ 869] = 1'b1; frame2.error[ 869] = 1'b0;frame2.data[ 870] = 8'h5B; frame2.valid[ 870] = 1'b1; frame2.error[ 870] = 1'b0;frame2.data[ 871] = 8'h5C; frame2.valid[ 871] = 1'b1; frame2.error[ 871] = 1'b0;frame2.data[ 872] = 8'h5D; frame2.valid[ 872] = 1'b1; frame2.error[ 872] = 1'b0;frame2.data[ 873] = 8'h5E; frame2.valid[ 873] = 1'b1; frame2.error[ 873] = 1'b0;frame2.data[ 874] = 8'h5F; frame2.valid[ 874] = 1'b1; frame2.error[ 874] = 1'b0;frame2.data[ 875] = 8'h60; frame2.valid[ 875] = 1'b1; frame2.error[ 875] = 1'b0;frame2.data[ 876] = 8'h61; frame2.valid[ 876] = 1'b1; frame2.error[ 876] = 1'b0;frame2.data[ 877] = 8'h62; frame2.valid[ 877] = 1'b1; frame2.error[ 877] = 1'b0;
        frame2.data[ 878] = 8'h63; frame2.valid[ 878] = 1'b1; frame2.error[ 878] = 1'b0;frame2.data[ 879] = 8'h64; frame2.valid[ 879] = 1'b1; frame2.error[ 879] = 1'b0;frame2.data[ 880] = 8'h65; frame2.valid[ 880] = 1'b1; frame2.error[ 880] = 1'b0;frame2.data[ 881] = 8'h66; frame2.valid[ 881] = 1'b1; frame2.error[ 881] = 1'b0;frame2.data[ 882] = 8'h67; frame2.valid[ 882] = 1'b1; frame2.error[ 882] = 1'b0;frame2.data[ 883] = 8'h68; frame2.valid[ 883] = 1'b1; frame2.error[ 883] = 1'b0;frame2.data[ 884] = 8'h69; frame2.valid[ 884] = 1'b1; frame2.error[ 884] = 1'b0;frame2.data[ 885] = 8'h6A; frame2.valid[ 885] = 1'b1; frame2.error[ 885] = 1'b0;frame2.data[ 886] = 8'h6B; frame2.valid[ 886] = 1'b1; frame2.error[ 886] = 1'b0;frame2.data[ 887] = 8'h6C; frame2.valid[ 887] = 1'b1; frame2.error[ 887] = 1'b0;frame2.data[ 888] = 8'h6D; frame2.valid[ 888] = 1'b1; frame2.error[ 888] = 1'b0;frame2.data[ 889] = 8'h6E; frame2.valid[ 889] = 1'b1; frame2.error[ 889] = 1'b0;frame2.data[ 890] = 8'h6F; frame2.valid[ 890] = 1'b1; frame2.error[ 890] = 1'b0;frame2.data[ 891] = 8'h70; frame2.valid[ 891] = 1'b1; frame2.error[ 891] = 1'b0;frame2.data[ 892] = 8'h71; frame2.valid[ 892] = 1'b1; frame2.error[ 892] = 1'b0;frame2.data[ 893] = 8'h72; frame2.valid[ 893] = 1'b1; frame2.error[ 893] = 1'b0;
        frame2.data[ 894] = 8'h73; frame2.valid[ 894] = 1'b1; frame2.error[ 894] = 1'b0;frame2.data[ 895] = 8'h74; frame2.valid[ 895] = 1'b1; frame2.error[ 895] = 1'b0;frame2.data[ 896] = 8'h75; frame2.valid[ 896] = 1'b1; frame2.error[ 896] = 1'b0;frame2.data[ 897] = 8'h76; frame2.valid[ 897] = 1'b1; frame2.error[ 897] = 1'b0;frame2.data[ 898] = 8'h77; frame2.valid[ 898] = 1'b1; frame2.error[ 898] = 1'b0;frame2.data[ 899] = 8'h78; frame2.valid[ 899] = 1'b1; frame2.error[ 899] = 1'b0;frame2.data[ 900] = 8'h79; frame2.valid[ 900] = 1'b1; frame2.error[ 900] = 1'b0;frame2.data[ 901] = 8'h7A; frame2.valid[ 901] = 1'b1; frame2.error[ 901] = 1'b0;frame2.data[ 902] = 8'h7B; frame2.valid[ 902] = 1'b1; frame2.error[ 902] = 1'b0;frame2.data[ 903] = 8'h7C; frame2.valid[ 903] = 1'b1; frame2.error[ 903] = 1'b0;frame2.data[ 904] = 8'h7D; frame2.valid[ 904] = 1'b1; frame2.error[ 904] = 1'b0;frame2.data[ 905] = 8'h7E; frame2.valid[ 905] = 1'b1; frame2.error[ 905] = 1'b0;frame2.data[ 906] = 8'h7F; frame2.valid[ 906] = 1'b1; frame2.error[ 906] = 1'b0;frame2.data[ 907] = 8'h80; frame2.valid[ 907] = 1'b1; frame2.error[ 907] = 1'b0;frame2.data[ 908] = 8'h81; frame2.valid[ 908] = 1'b1; frame2.error[ 908] = 1'b0;frame2.data[ 909] = 8'h82; frame2.valid[ 909] = 1'b1; frame2.error[ 909] = 1'b0;
        frame2.data[ 910] = 8'h83; frame2.valid[ 910] = 1'b1; frame2.error[ 910] = 1'b0;frame2.data[ 911] = 8'h84; frame2.valid[ 911] = 1'b1; frame2.error[ 911] = 1'b0;frame2.data[ 912] = 8'h85; frame2.valid[ 912] = 1'b1; frame2.error[ 912] = 1'b0;frame2.data[ 913] = 8'h86; frame2.valid[ 913] = 1'b1; frame2.error[ 913] = 1'b0;frame2.data[ 914] = 8'h87; frame2.valid[ 914] = 1'b1; frame2.error[ 914] = 1'b0;frame2.data[ 915] = 8'h88; frame2.valid[ 915] = 1'b1; frame2.error[ 915] = 1'b0;frame2.data[ 916] = 8'h89; frame2.valid[ 916] = 1'b1; frame2.error[ 916] = 1'b0;frame2.data[ 917] = 8'h8A; frame2.valid[ 917] = 1'b1; frame2.error[ 917] = 1'b0;frame2.data[ 918] = 8'h8B; frame2.valid[ 918] = 1'b1; frame2.error[ 918] = 1'b0;frame2.data[ 919] = 8'h8C; frame2.valid[ 919] = 1'b1; frame2.error[ 919] = 1'b0;frame2.data[ 920] = 8'h8D; frame2.valid[ 920] = 1'b1; frame2.error[ 920] = 1'b0;frame2.data[ 921] = 8'h8E; frame2.valid[ 921] = 1'b1; frame2.error[ 921] = 1'b0;frame2.data[ 922] = 8'h8F; frame2.valid[ 922] = 1'b1; frame2.error[ 922] = 1'b0;frame2.data[ 923] = 8'h90; frame2.valid[ 923] = 1'b1; frame2.error[ 923] = 1'b0;frame2.data[ 924] = 8'h91; frame2.valid[ 924] = 1'b1; frame2.error[ 924] = 1'b0;frame2.data[ 925] = 8'h92; frame2.valid[ 925] = 1'b1; frame2.error[ 925] = 1'b0;
        frame2.data[ 926] = 8'h93; frame2.valid[ 926] = 1'b1; frame2.error[ 926] = 1'b0;frame2.data[ 927] = 8'h94; frame2.valid[ 927] = 1'b1; frame2.error[ 927] = 1'b0;frame2.data[ 928] = 8'h95; frame2.valid[ 928] = 1'b1; frame2.error[ 928] = 1'b0;frame2.data[ 929] = 8'h96; frame2.valid[ 929] = 1'b1; frame2.error[ 929] = 1'b0;frame2.data[ 930] = 8'h97; frame2.valid[ 930] = 1'b1; frame2.error[ 930] = 1'b0;frame2.data[ 931] = 8'h98; frame2.valid[ 931] = 1'b1; frame2.error[ 931] = 1'b0;frame2.data[ 932] = 8'h99; frame2.valid[ 932] = 1'b1; frame2.error[ 932] = 1'b0;frame2.data[ 933] = 8'h9A; frame2.valid[ 933] = 1'b1; frame2.error[ 933] = 1'b0;frame2.data[ 934] = 8'h9B; frame2.valid[ 934] = 1'b1; frame2.error[ 934] = 1'b0;frame2.data[ 935] = 8'h9C; frame2.valid[ 935] = 1'b1; frame2.error[ 935] = 1'b0;frame2.data[ 936] = 8'h9D; frame2.valid[ 936] = 1'b1; frame2.error[ 936] = 1'b0;frame2.data[ 937] = 8'h9E; frame2.valid[ 937] = 1'b1; frame2.error[ 937] = 1'b0;frame2.data[ 938] = 8'h9F; frame2.valid[ 938] = 1'b1; frame2.error[ 938] = 1'b0;frame2.data[ 939] = 8'hA0; frame2.valid[ 939] = 1'b1; frame2.error[ 939] = 1'b0;frame2.data[ 940] = 8'hA1; frame2.valid[ 940] = 1'b1; frame2.error[ 940] = 1'b0;frame2.data[ 941] = 8'hA2; frame2.valid[ 941] = 1'b1; frame2.error[ 941] = 1'b0;
        frame2.data[ 942] = 8'hA3; frame2.valid[ 942] = 1'b1; frame2.error[ 942] = 1'b0;frame2.data[ 943] = 8'hA4; frame2.valid[ 943] = 1'b1; frame2.error[ 943] = 1'b0;frame2.data[ 944] = 8'hA5; frame2.valid[ 944] = 1'b1; frame2.error[ 944] = 1'b0;frame2.data[ 945] = 8'hA6; frame2.valid[ 945] = 1'b1; frame2.error[ 945] = 1'b0;frame2.data[ 946] = 8'hA7; frame2.valid[ 946] = 1'b1; frame2.error[ 946] = 1'b0;frame2.data[ 947] = 8'hA8; frame2.valid[ 947] = 1'b1; frame2.error[ 947] = 1'b0;frame2.data[ 948] = 8'hA9; frame2.valid[ 948] = 1'b1; frame2.error[ 948] = 1'b0;frame2.data[ 949] = 8'hAA; frame2.valid[ 949] = 1'b1; frame2.error[ 949] = 1'b0;frame2.data[ 950] = 8'hAB; frame2.valid[ 950] = 1'b1; frame2.error[ 950] = 1'b0;frame2.data[ 951] = 8'hAC; frame2.valid[ 951] = 1'b1; frame2.error[ 951] = 1'b0;frame2.data[ 952] = 8'hAD; frame2.valid[ 952] = 1'b1; frame2.error[ 952] = 1'b0;frame2.data[ 953] = 8'hAE; frame2.valid[ 953] = 1'b1; frame2.error[ 953] = 1'b0;frame2.data[ 954] = 8'hAF; frame2.valid[ 954] = 1'b1; frame2.error[ 954] = 1'b0;frame2.data[ 955] = 8'hB0; frame2.valid[ 955] = 1'b1; frame2.error[ 955] = 1'b0;frame2.data[ 956] = 8'hB1; frame2.valid[ 956] = 1'b1; frame2.error[ 956] = 1'b0;frame2.data[ 957] = 8'hB2; frame2.valid[ 957] = 1'b1; frame2.error[ 957] = 1'b0;
        frame2.data[ 958] = 8'hB3; frame2.valid[ 958] = 1'b1; frame2.error[ 958] = 1'b0;frame2.data[ 959] = 8'hB4; frame2.valid[ 959] = 1'b1; frame2.error[ 959] = 1'b0;frame2.data[ 960] = 8'hB5; frame2.valid[ 960] = 1'b1; frame2.error[ 960] = 1'b0;frame2.data[ 961] = 8'hB6; frame2.valid[ 961] = 1'b1; frame2.error[ 961] = 1'b0;frame2.data[ 962] = 8'hB7; frame2.valid[ 962] = 1'b1; frame2.error[ 962] = 1'b0;frame2.data[ 963] = 8'hB8; frame2.valid[ 963] = 1'b1; frame2.error[ 963] = 1'b0;frame2.data[ 964] = 8'hB9; frame2.valid[ 964] = 1'b1; frame2.error[ 964] = 1'b0;frame2.data[ 965] = 8'hBA; frame2.valid[ 965] = 1'b1; frame2.error[ 965] = 1'b0;frame2.data[ 966] = 8'hBB; frame2.valid[ 966] = 1'b1; frame2.error[ 966] = 1'b0;frame2.data[ 967] = 8'hBC; frame2.valid[ 967] = 1'b1; frame2.error[ 967] = 1'b0;frame2.data[ 968] = 8'hBD; frame2.valid[ 968] = 1'b1; frame2.error[ 968] = 1'b0;frame2.data[ 969] = 8'hBE; frame2.valid[ 969] = 1'b1; frame2.error[ 969] = 1'b0;frame2.data[ 970] = 8'hBF; frame2.valid[ 970] = 1'b1; frame2.error[ 970] = 1'b0;frame2.data[ 971] = 8'hC0; frame2.valid[ 971] = 1'b1; frame2.error[ 971] = 1'b0;frame2.data[ 972] = 8'hC1; frame2.valid[ 972] = 1'b1; frame2.error[ 972] = 1'b0;frame2.data[ 973] = 8'hC2; frame2.valid[ 973] = 1'b1; frame2.error[ 973] = 1'b0;
        frame2.data[ 974] = 8'hC3; frame2.valid[ 974] = 1'b1; frame2.error[ 974] = 1'b0;frame2.data[ 975] = 8'hC4; frame2.valid[ 975] = 1'b1; frame2.error[ 975] = 1'b0;frame2.data[ 976] = 8'hC5; frame2.valid[ 976] = 1'b1; frame2.error[ 976] = 1'b0;frame2.data[ 977] = 8'hC6; frame2.valid[ 977] = 1'b1; frame2.error[ 977] = 1'b0;frame2.data[ 978] = 8'hC7; frame2.valid[ 978] = 1'b1; frame2.error[ 978] = 1'b0;frame2.data[ 979] = 8'hC8; frame2.valid[ 979] = 1'b1; frame2.error[ 979] = 1'b0;frame2.data[ 980] = 8'hC9; frame2.valid[ 980] = 1'b1; frame2.error[ 980] = 1'b0;frame2.data[ 981] = 8'hCA; frame2.valid[ 981] = 1'b1; frame2.error[ 981] = 1'b0;frame2.data[ 982] = 8'hCB; frame2.valid[ 982] = 1'b1; frame2.error[ 982] = 1'b0;frame2.data[ 983] = 8'hCC; frame2.valid[ 983] = 1'b1; frame2.error[ 983] = 1'b0;frame2.data[ 984] = 8'hCD; frame2.valid[ 984] = 1'b1; frame2.error[ 984] = 1'b0;frame2.data[ 985] = 8'hCE; frame2.valid[ 985] = 1'b1; frame2.error[ 985] = 1'b0;frame2.data[ 986] = 8'hCF; frame2.valid[ 986] = 1'b1; frame2.error[ 986] = 1'b0;frame2.data[ 987] = 8'hD0; frame2.valid[ 987] = 1'b1; frame2.error[ 987] = 1'b0;frame2.data[ 988] = 8'hD1; frame2.valid[ 988] = 1'b1; frame2.error[ 988] = 1'b0;frame2.data[ 989] = 8'hD2; frame2.valid[ 989] = 1'b1; frame2.error[ 989] = 1'b0;
        frame2.data[ 990] = 8'hD3; frame2.valid[ 990] = 1'b1; frame2.error[ 990] = 1'b0;frame2.data[ 991] = 8'hD4; frame2.valid[ 991] = 1'b1; frame2.error[ 991] = 1'b0;frame2.data[ 992] = 8'hD5; frame2.valid[ 992] = 1'b1; frame2.error[ 992] = 1'b0;frame2.data[ 993] = 8'hD6; frame2.valid[ 993] = 1'b1; frame2.error[ 993] = 1'b0;frame2.data[ 994] = 8'hD7; frame2.valid[ 994] = 1'b1; frame2.error[ 994] = 1'b0;frame2.data[ 995] = 8'hD8; frame2.valid[ 995] = 1'b1; frame2.error[ 995] = 1'b0;frame2.data[ 996] = 8'hD9; frame2.valid[ 996] = 1'b1; frame2.error[ 996] = 1'b0;frame2.data[ 997] = 8'hDA; frame2.valid[ 997] = 1'b1; frame2.error[ 997] = 1'b0;frame2.data[ 998] = 8'hDB; frame2.valid[ 998] = 1'b1; frame2.error[ 998] = 1'b0;frame2.data[ 999] = 8'hDC; frame2.valid[ 999] = 1'b1; frame2.error[ 999] = 1'b0;frame2.data[1000] = 8'hDD; frame2.valid[1000] = 1'b1; frame2.error[1000] = 1'b0;frame2.data[1001] = 8'hDE; frame2.valid[1001] = 1'b1; frame2.error[1001] = 1'b0;frame2.data[1002] = 8'hDF; frame2.valid[1002] = 1'b1; frame2.error[1002] = 1'b0;frame2.data[1003] = 8'hE0; frame2.valid[1003] = 1'b1; frame2.error[1003] = 1'b0;frame2.data[1004] = 8'hE1; frame2.valid[1004] = 1'b1; frame2.error[1004] = 1'b0;frame2.data[1005] = 8'hE2; frame2.valid[1005] = 1'b1; frame2.error[1005] = 1'b0;
        frame2.data[1006] = 8'hE3; frame2.valid[1006] = 1'b1; frame2.error[1006] = 1'b0;frame2.data[1007] = 8'hE4; frame2.valid[1007] = 1'b1; frame2.error[1007] = 1'b0;frame2.data[1008] = 8'hE5; frame2.valid[1008] = 1'b1; frame2.error[1008] = 1'b0;frame2.data[1009] = 8'hE6; frame2.valid[1009] = 1'b1; frame2.error[1009] = 1'b0;frame2.data[1010] = 8'hE7; frame2.valid[1010] = 1'b1; frame2.error[1010] = 1'b0;frame2.data[1011] = 8'hE8; frame2.valid[1011] = 1'b1; frame2.error[1011] = 1'b0;frame2.data[1012] = 8'hE9; frame2.valid[1012] = 1'b1; frame2.error[1012] = 1'b0;frame2.data[1013] = 8'hEA; frame2.valid[1013] = 1'b1; frame2.error[1013] = 1'b0;frame2.data[1014] = 8'hEB; frame2.valid[1014] = 1'b1; frame2.error[1014] = 1'b0;frame2.data[1015] = 8'hEC; frame2.valid[1015] = 1'b1; frame2.error[1015] = 1'b0;frame2.data[1016] = 8'hED; frame2.valid[1016] = 1'b1; frame2.error[1016] = 1'b0;frame2.data[1017] = 8'hEE; frame2.valid[1017] = 1'b1; frame2.error[1017] = 1'b0;frame2.data[1018] = 8'hEF; frame2.valid[1018] = 1'b1; frame2.error[1018] = 1'b0;frame2.data[1019] = 8'hF0; frame2.valid[1019] = 1'b1; frame2.error[1019] = 1'b0;frame2.data[1020] = 8'hF1; frame2.valid[1020] = 1'b1; frame2.error[1020] = 1'b0;frame2.data[1021] = 8'hF2; frame2.valid[1021] = 1'b1; frame2.error[1021] = 1'b0;
        frame2.data[1022] = 8'hF3; frame2.valid[1022] = 1'b1; frame2.error[1022] = 1'b0;frame2.data[1023] = 8'hF4; frame2.valid[1023] = 1'b1; frame2.error[1023] = 1'b0;frame2.data[1024] = 8'hF5; frame2.valid[1024] = 1'b1; frame2.error[1024] = 1'b0;frame2.data[1025] = 8'hF6; frame2.valid[1025] = 1'b1; frame2.error[1025] = 1'b0;frame2.data[1026] = 8'hF7; frame2.valid[1026] = 1'b1; frame2.error[1026] = 1'b0;frame2.data[1027] = 8'hF8; frame2.valid[1027] = 1'b1; frame2.error[1027] = 1'b0;frame2.data[1028] = 8'hF9; frame2.valid[1028] = 1'b1; frame2.error[1028] = 1'b0;frame2.data[1029] = 8'hFA; frame2.valid[1029] = 1'b1; frame2.error[1029] = 1'b0;frame2.data[1030] = 8'hFB; frame2.valid[1030] = 1'b1; frame2.error[1030] = 1'b0;frame2.data[1031] = 8'hFC; frame2.valid[1031] = 1'b1; frame2.error[1031] = 1'b0;frame2.data[1032] = 8'hFD; frame2.valid[1032] = 1'b1; frame2.error[1032] = 1'b0;frame2.data[1033] = 8'hFE; frame2.valid[1033] = 1'b1; frame2.error[1033] = 1'b0;frame2.data[1034] = 8'h00; frame2.valid[1034] = 1'b1; frame2.error[1034] = 1'b0;frame2.data[1035] = 8'h01; frame2.valid[1035] = 1'b1; frame2.error[1035] = 1'b0;frame2.data[1036] = 8'h02; frame2.valid[1036] = 1'b1; frame2.error[1036] = 1'b0;frame2.data[1037] = 8'h03; frame2.valid[1037] = 1'b1; frame2.error[1037] = 1'b0;
        frame2.data[1038] = 8'h04; frame2.valid[1038] = 1'b1; frame2.error[1038] = 1'b0;frame2.data[1039] = 8'h05; frame2.valid[1039] = 1'b1; frame2.error[1039] = 1'b0;frame2.data[1040] = 8'h06; frame2.valid[1040] = 1'b1; frame2.error[1040] = 1'b0;frame2.data[1041] = 8'h07; frame2.valid[1041] = 1'b1; frame2.error[1041] = 1'b0;frame2.data[1042] = 8'h08; frame2.valid[1042] = 1'b1; frame2.error[1042] = 1'b0;frame2.data[1043] = 8'h09; frame2.valid[1043] = 1'b1; frame2.error[1043] = 1'b0;frame2.data[1044] = 8'h0A; frame2.valid[1044] = 1'b1; frame2.error[1044] = 1'b0;frame2.data[1045] = 8'h0B; frame2.valid[1045] = 1'b1; frame2.error[1045] = 1'b0;frame2.data[1046] = 8'h0C; frame2.valid[1046] = 1'b1; frame2.error[1046] = 1'b0;frame2.data[1047] = 8'h0D; frame2.valid[1047] = 1'b1; frame2.error[1047] = 1'b0;frame2.data[1048] = 8'h0E; frame2.valid[1048] = 1'b1; frame2.error[1048] = 1'b0;frame2.data[1049] = 8'h0F; frame2.valid[1049] = 1'b1; frame2.error[1049] = 1'b0;frame2.data[1050] = 8'h10; frame2.valid[1050] = 1'b1; frame2.error[1050] = 1'b0;frame2.data[1051] = 8'h11; frame2.valid[1051] = 1'b1; frame2.error[1051] = 1'b0;frame2.data[1052] = 8'h12; frame2.valid[1052] = 1'b1; frame2.error[1052] = 1'b0;frame2.data[1053] = 8'h13; frame2.valid[1053] = 1'b1; frame2.error[1053] = 1'b0;
        frame2.data[1054] = 8'h14; frame2.valid[1054] = 1'b1; frame2.error[1054] = 1'b0;frame2.data[1055] = 8'h15; frame2.valid[1055] = 1'b1; frame2.error[1055] = 1'b0;frame2.data[1056] = 8'h16; frame2.valid[1056] = 1'b1; frame2.error[1056] = 1'b0;frame2.data[1057] = 8'h17; frame2.valid[1057] = 1'b1; frame2.error[1057] = 1'b0;frame2.data[1058] = 8'h18; frame2.valid[1058] = 1'b1; frame2.error[1058] = 1'b0;frame2.data[1059] = 8'h19; frame2.valid[1059] = 1'b1; frame2.error[1059] = 1'b0;frame2.data[1060] = 8'h1A; frame2.valid[1060] = 1'b1; frame2.error[1060] = 1'b0;frame2.data[1061] = 8'h1B; frame2.valid[1061] = 1'b1; frame2.error[1061] = 1'b0;frame2.data[1062] = 8'h1C; frame2.valid[1062] = 1'b1; frame2.error[1062] = 1'b0;frame2.data[1063] = 8'h1D; frame2.valid[1063] = 1'b1; frame2.error[1063] = 1'b0;frame2.data[1064] = 8'h1E; frame2.valid[1064] = 1'b1; frame2.error[1064] = 1'b0;frame2.data[1065] = 8'h1F; frame2.valid[1065] = 1'b1; frame2.error[1065] = 1'b0;frame2.data[1066] = 8'h20; frame2.valid[1066] = 1'b1; frame2.error[1066] = 1'b0;frame2.data[1067] = 8'h21; frame2.valid[1067] = 1'b1; frame2.error[1067] = 1'b0;frame2.data[1068] = 8'h22; frame2.valid[1068] = 1'b1; frame2.error[1068] = 1'b0;frame2.data[1069] = 8'h23; frame2.valid[1069] = 1'b1; frame2.error[1069] = 1'b0;
        frame2.data[1070] = 8'h24; frame2.valid[1070] = 1'b1; frame2.error[1070] = 1'b0;frame2.data[1071] = 8'h25; frame2.valid[1071] = 1'b1; frame2.error[1071] = 1'b0;frame2.data[1072] = 8'h26; frame2.valid[1072] = 1'b1; frame2.error[1072] = 1'b0;frame2.data[1073] = 8'h27; frame2.valid[1073] = 1'b1; frame2.error[1073] = 1'b0;frame2.data[1074] = 8'h28; frame2.valid[1074] = 1'b1; frame2.error[1074] = 1'b0;frame2.data[1075] = 8'h29; frame2.valid[1075] = 1'b1; frame2.error[1075] = 1'b0;frame2.data[1076] = 8'h2A; frame2.valid[1076] = 1'b1; frame2.error[1076] = 1'b0;frame2.data[1077] = 8'h2B; frame2.valid[1077] = 1'b1; frame2.error[1077] = 1'b0;frame2.data[1078] = 8'h2C; frame2.valid[1078] = 1'b1; frame2.error[1078] = 1'b0;frame2.data[1079] = 8'h2D; frame2.valid[1079] = 1'b1; frame2.error[1079] = 1'b0;frame2.data[1080] = 8'h2E; frame2.valid[1080] = 1'b1; frame2.error[1080] = 1'b0;frame2.data[1081] = 8'h2F; frame2.valid[1081] = 1'b1; frame2.error[1081] = 1'b0;frame2.data[1082] = 8'h30; frame2.valid[1082] = 1'b1; frame2.error[1082] = 1'b0;frame2.data[1083] = 8'h31; frame2.valid[1083] = 1'b1; frame2.error[1083] = 1'b0;frame2.data[1084] = 8'h32; frame2.valid[1084] = 1'b1; frame2.error[1084] = 1'b0;frame2.data[1085] = 8'h33; frame2.valid[1085] = 1'b1; frame2.error[1085] = 1'b0;
        frame2.data[1086] = 8'h34; frame2.valid[1086] = 1'b1; frame2.error[1086] = 1'b0;frame2.data[1087] = 8'h35; frame2.valid[1087] = 1'b1; frame2.error[1087] = 1'b0;frame2.data[1088] = 8'h36; frame2.valid[1088] = 1'b1; frame2.error[1088] = 1'b0;frame2.data[1089] = 8'h37; frame2.valid[1089] = 1'b1; frame2.error[1089] = 1'b0;frame2.data[1090] = 8'h38; frame2.valid[1090] = 1'b1; frame2.error[1090] = 1'b0;frame2.data[1091] = 8'h39; frame2.valid[1091] = 1'b1; frame2.error[1091] = 1'b0;frame2.data[1092] = 8'h3A; frame2.valid[1092] = 1'b1; frame2.error[1092] = 1'b0;frame2.data[1093] = 8'h3B; frame2.valid[1093] = 1'b1; frame2.error[1093] = 1'b0;frame2.data[1094] = 8'h3C; frame2.valid[1094] = 1'b1; frame2.error[1094] = 1'b0;frame2.data[1095] = 8'h3D; frame2.valid[1095] = 1'b1; frame2.error[1095] = 1'b0;frame2.data[1096] = 8'h3E; frame2.valid[1096] = 1'b1; frame2.error[1096] = 1'b0;frame2.data[1097] = 8'h3F; frame2.valid[1097] = 1'b1; frame2.error[1097] = 1'b0;frame2.data[1098] = 8'h40; frame2.valid[1098] = 1'b1; frame2.error[1098] = 1'b0;frame2.data[1099] = 8'h41; frame2.valid[1099] = 1'b1; frame2.error[1099] = 1'b0;frame2.data[1100] = 8'h42; frame2.valid[1100] = 1'b1; frame2.error[1100] = 1'b0;frame2.data[1101] = 8'h43; frame2.valid[1101] = 1'b1; frame2.error[1101] = 1'b0;
        frame2.data[1102] = 8'h44; frame2.valid[1102] = 1'b1; frame2.error[1102] = 1'b0;frame2.data[1103] = 8'h45; frame2.valid[1103] = 1'b1; frame2.error[1103] = 1'b0;frame2.data[1104] = 8'h46; frame2.valid[1104] = 1'b1; frame2.error[1104] = 1'b0;frame2.data[1105] = 8'h47; frame2.valid[1105] = 1'b1; frame2.error[1105] = 1'b0;frame2.data[1106] = 8'h48; frame2.valid[1106] = 1'b1; frame2.error[1106] = 1'b0;frame2.data[1107] = 8'h49; frame2.valid[1107] = 1'b1; frame2.error[1107] = 1'b0;frame2.data[1108] = 8'h4A; frame2.valid[1108] = 1'b1; frame2.error[1108] = 1'b0;frame2.data[1109] = 8'h4B; frame2.valid[1109] = 1'b1; frame2.error[1109] = 1'b0;frame2.data[1110] = 8'h4C; frame2.valid[1110] = 1'b1; frame2.error[1110] = 1'b0;frame2.data[1111] = 8'h4D; frame2.valid[1111] = 1'b1; frame2.error[1111] = 1'b0;frame2.data[1112] = 8'h4E; frame2.valid[1112] = 1'b1; frame2.error[1112] = 1'b0;frame2.data[1113] = 8'h4F; frame2.valid[1113] = 1'b1; frame2.error[1113] = 1'b0;frame2.data[1114] = 8'h50; frame2.valid[1114] = 1'b1; frame2.error[1114] = 1'b0;frame2.data[1115] = 8'h51; frame2.valid[1115] = 1'b1; frame2.error[1115] = 1'b0;frame2.data[1116] = 8'h52; frame2.valid[1116] = 1'b1; frame2.error[1116] = 1'b0;frame2.data[1117] = 8'h53; frame2.valid[1117] = 1'b1; frame2.error[1117] = 1'b0;
        frame2.data[1118] = 8'h54; frame2.valid[1118] = 1'b1; frame2.error[1118] = 1'b0;frame2.data[1119] = 8'h55; frame2.valid[1119] = 1'b1; frame2.error[1119] = 1'b0;frame2.data[1120] = 8'h56; frame2.valid[1120] = 1'b1; frame2.error[1120] = 1'b0;frame2.data[1121] = 8'h57; frame2.valid[1121] = 1'b1; frame2.error[1121] = 1'b0;frame2.data[1122] = 8'h58; frame2.valid[1122] = 1'b1; frame2.error[1122] = 1'b0;frame2.data[1123] = 8'h59; frame2.valid[1123] = 1'b1; frame2.error[1123] = 1'b0;frame2.data[1124] = 8'h5A; frame2.valid[1124] = 1'b1; frame2.error[1124] = 1'b0;frame2.data[1125] = 8'h5B; frame2.valid[1125] = 1'b1; frame2.error[1125] = 1'b0;frame2.data[1126] = 8'h5C; frame2.valid[1126] = 1'b1; frame2.error[1126] = 1'b0;frame2.data[1127] = 8'h5D; frame2.valid[1127] = 1'b1; frame2.error[1127] = 1'b0;frame2.data[1128] = 8'h5E; frame2.valid[1128] = 1'b1; frame2.error[1128] = 1'b0;frame2.data[1129] = 8'h5F; frame2.valid[1129] = 1'b1; frame2.error[1129] = 1'b0;frame2.data[1130] = 8'h60; frame2.valid[1130] = 1'b1; frame2.error[1130] = 1'b0;frame2.data[1131] = 8'h61; frame2.valid[1131] = 1'b1; frame2.error[1131] = 1'b0;frame2.data[1132] = 8'h62; frame2.valid[1132] = 1'b1; frame2.error[1132] = 1'b0;frame2.data[1133] = 8'h63; frame2.valid[1133] = 1'b1; frame2.error[1133] = 1'b0;
        frame2.data[1134] = 8'h64; frame2.valid[1134] = 1'b1; frame2.error[1134] = 1'b0;frame2.data[1135] = 8'h65; frame2.valid[1135] = 1'b1; frame2.error[1135] = 1'b0;frame2.data[1136] = 8'h66; frame2.valid[1136] = 1'b1; frame2.error[1136] = 1'b0;frame2.data[1137] = 8'h67; frame2.valid[1137] = 1'b1; frame2.error[1137] = 1'b0;frame2.data[1138] = 8'h68; frame2.valid[1138] = 1'b1; frame2.error[1138] = 1'b0;frame2.data[1139] = 8'h69; frame2.valid[1139] = 1'b1; frame2.error[1139] = 1'b0;frame2.data[1140] = 8'h6A; frame2.valid[1140] = 1'b1; frame2.error[1140] = 1'b0;frame2.data[1141] = 8'h6B; frame2.valid[1141] = 1'b1; frame2.error[1141] = 1'b0;frame2.data[1142] = 8'h6C; frame2.valid[1142] = 1'b1; frame2.error[1142] = 1'b0;frame2.data[1143] = 8'h6D; frame2.valid[1143] = 1'b1; frame2.error[1143] = 1'b0;frame2.data[1144] = 8'h6E; frame2.valid[1144] = 1'b1; frame2.error[1144] = 1'b0;frame2.data[1145] = 8'h6F; frame2.valid[1145] = 1'b1; frame2.error[1145] = 1'b0;frame2.data[1146] = 8'h70; frame2.valid[1146] = 1'b1; frame2.error[1146] = 1'b0;frame2.data[1147] = 8'h71; frame2.valid[1147] = 1'b1; frame2.error[1147] = 1'b0;frame2.data[1148] = 8'h72; frame2.valid[1148] = 1'b1; frame2.error[1148] = 1'b0;frame2.data[1149] = 8'h73; frame2.valid[1149] = 1'b1; frame2.error[1149] = 1'b0;
        frame2.data[1150] = 8'h74; frame2.valid[1150] = 1'b1; frame2.error[1150] = 1'b0;frame2.data[1151] = 8'h75; frame2.valid[1151] = 1'b1; frame2.error[1151] = 1'b0;frame2.data[1152] = 8'h76; frame2.valid[1152] = 1'b1; frame2.error[1152] = 1'b0;frame2.data[1153] = 8'h77; frame2.valid[1153] = 1'b1; frame2.error[1153] = 1'b0;frame2.data[1154] = 8'h78; frame2.valid[1154] = 1'b1; frame2.error[1154] = 1'b0;frame2.data[1155] = 8'h79; frame2.valid[1155] = 1'b1; frame2.error[1155] = 1'b0;frame2.data[1156] = 8'h7A; frame2.valid[1156] = 1'b1; frame2.error[1156] = 1'b0;frame2.data[1157] = 8'h7B; frame2.valid[1157] = 1'b1; frame2.error[1157] = 1'b0;frame2.data[1158] = 8'h7C; frame2.valid[1158] = 1'b1; frame2.error[1158] = 1'b0;frame2.data[1159] = 8'h7D; frame2.valid[1159] = 1'b1; frame2.error[1159] = 1'b0;frame2.data[1160] = 8'h7E; frame2.valid[1160] = 1'b1; frame2.error[1160] = 1'b0;frame2.data[1161] = 8'h7F; frame2.valid[1161] = 1'b1; frame2.error[1161] = 1'b0;frame2.data[1162] = 8'h80; frame2.valid[1162] = 1'b1; frame2.error[1162] = 1'b0;frame2.data[1163] = 8'h81; frame2.valid[1163] = 1'b1; frame2.error[1163] = 1'b0;frame2.data[1164] = 8'h82; frame2.valid[1164] = 1'b1; frame2.error[1164] = 1'b0;frame2.data[1165] = 8'h83; frame2.valid[1165] = 1'b1; frame2.error[1165] = 1'b0;
        frame2.data[1166] = 8'h84; frame2.valid[1166] = 1'b1; frame2.error[1166] = 1'b0;frame2.data[1167] = 8'h85; frame2.valid[1167] = 1'b1; frame2.error[1167] = 1'b0;frame2.data[1168] = 8'h86; frame2.valid[1168] = 1'b1; frame2.error[1168] = 1'b0;frame2.data[1169] = 8'h87; frame2.valid[1169] = 1'b1; frame2.error[1169] = 1'b0;frame2.data[1170] = 8'h88; frame2.valid[1170] = 1'b1; frame2.error[1170] = 1'b0;frame2.data[1171] = 8'h89; frame2.valid[1171] = 1'b1; frame2.error[1171] = 1'b0;frame2.data[1172] = 8'h8A; frame2.valid[1172] = 1'b1; frame2.error[1172] = 1'b0;frame2.data[1173] = 8'h8B; frame2.valid[1173] = 1'b1; frame2.error[1173] = 1'b0;frame2.data[1174] = 8'h8C; frame2.valid[1174] = 1'b1; frame2.error[1174] = 1'b0;frame2.data[1175] = 8'h8D; frame2.valid[1175] = 1'b1; frame2.error[1175] = 1'b0;frame2.data[1176] = 8'h8E; frame2.valid[1176] = 1'b1; frame2.error[1176] = 1'b0;frame2.data[1177] = 8'h8F; frame2.valid[1177] = 1'b1; frame2.error[1177] = 1'b0;frame2.data[1178] = 8'h90; frame2.valid[1178] = 1'b1; frame2.error[1178] = 1'b0;frame2.data[1179] = 8'h91; frame2.valid[1179] = 1'b1; frame2.error[1179] = 1'b0;frame2.data[1180] = 8'h92; frame2.valid[1180] = 1'b1; frame2.error[1180] = 1'b0;frame2.data[1181] = 8'h93; frame2.valid[1181] = 1'b1; frame2.error[1181] = 1'b0;
        frame2.data[1182] = 8'h94; frame2.valid[1182] = 1'b1; frame2.error[1182] = 1'b0;frame2.data[1183] = 8'h95; frame2.valid[1183] = 1'b1; frame2.error[1183] = 1'b0;frame2.data[1184] = 8'h96; frame2.valid[1184] = 1'b1; frame2.error[1184] = 1'b0;frame2.data[1185] = 8'h97; frame2.valid[1185] = 1'b1; frame2.error[1185] = 1'b0;frame2.data[1186] = 8'h98; frame2.valid[1186] = 1'b1; frame2.error[1186] = 1'b0;frame2.data[1187] = 8'h99; frame2.valid[1187] = 1'b1; frame2.error[1187] = 1'b0;frame2.data[1188] = 8'h9A; frame2.valid[1188] = 1'b1; frame2.error[1188] = 1'b0;frame2.data[1189] = 8'h9B; frame2.valid[1189] = 1'b1; frame2.error[1189] = 1'b0;frame2.data[1190] = 8'h9C; frame2.valid[1190] = 1'b1; frame2.error[1190] = 1'b0;frame2.data[1191] = 8'h9D; frame2.valid[1191] = 1'b1; frame2.error[1191] = 1'b0;frame2.data[1192] = 8'h9E; frame2.valid[1192] = 1'b1; frame2.error[1192] = 1'b0;frame2.data[1193] = 8'h9F; frame2.valid[1193] = 1'b1; frame2.error[1193] = 1'b0;frame2.data[1194] = 8'hA0; frame2.valid[1194] = 1'b1; frame2.error[1194] = 1'b0;frame2.data[1195] = 8'hA1; frame2.valid[1195] = 1'b1; frame2.error[1195] = 1'b0;frame2.data[1196] = 8'hA2; frame2.valid[1196] = 1'b1; frame2.error[1196] = 1'b0;frame2.data[1197] = 8'hA3; frame2.valid[1197] = 1'b1; frame2.error[1197] = 1'b0;
        frame2.data[1198] = 8'hA4; frame2.valid[1198] = 1'b1; frame2.error[1198] = 1'b0;frame2.data[1199] = 8'hA5; frame2.valid[1199] = 1'b1; frame2.error[1199] = 1'b0;frame2.data[1200] = 8'hA6; frame2.valid[1200] = 1'b1; frame2.error[1200] = 1'b0;frame2.data[1201] = 8'hA7; frame2.valid[1201] = 1'b1; frame2.error[1201] = 1'b0;frame2.data[1202] = 8'hA8; frame2.valid[1202] = 1'b1; frame2.error[1202] = 1'b0;frame2.data[1203] = 8'hA9; frame2.valid[1203] = 1'b1; frame2.error[1203] = 1'b0;frame2.data[1204] = 8'hAA; frame2.valid[1204] = 1'b1; frame2.error[1204] = 1'b0;frame2.data[1205] = 8'hAB; frame2.valid[1205] = 1'b1; frame2.error[1205] = 1'b0;frame2.data[1206] = 8'hAC; frame2.valid[1206] = 1'b1; frame2.error[1206] = 1'b0;frame2.data[1207] = 8'hAD; frame2.valid[1207] = 1'b1; frame2.error[1207] = 1'b0;frame2.data[1208] = 8'hAE; frame2.valid[1208] = 1'b1; frame2.error[1208] = 1'b0;frame2.data[1209] = 8'hAF; frame2.valid[1209] = 1'b1; frame2.error[1209] = 1'b0;frame2.data[1210] = 8'hB0; frame2.valid[1210] = 1'b1; frame2.error[1210] = 1'b0;frame2.data[1211] = 8'hB1; frame2.valid[1211] = 1'b1; frame2.error[1211] = 1'b0;frame2.data[1212] = 8'hB2; frame2.valid[1212] = 1'b1; frame2.error[1212] = 1'b0;frame2.data[1213] = 8'hB3; frame2.valid[1213] = 1'b1; frame2.error[1213] = 1'b0;
        frame2.data[1214] = 8'hB4; frame2.valid[1214] = 1'b1; frame2.error[1214] = 1'b0;frame2.data[1215] = 8'hB5; frame2.valid[1215] = 1'b1; frame2.error[1215] = 1'b0;frame2.data[1216] = 8'hB6; frame2.valid[1216] = 1'b1; frame2.error[1216] = 1'b0;frame2.data[1217] = 8'hB7; frame2.valid[1217] = 1'b1; frame2.error[1217] = 1'b0;frame2.data[1218] = 8'hB8; frame2.valid[1218] = 1'b1; frame2.error[1218] = 1'b0;frame2.data[1219] = 8'hB9; frame2.valid[1219] = 1'b1; frame2.error[1219] = 1'b0;frame2.data[1220] = 8'hBA; frame2.valid[1220] = 1'b1; frame2.error[1220] = 1'b0;frame2.data[1221] = 8'hBB; frame2.valid[1221] = 1'b1; frame2.error[1221] = 1'b0;frame2.data[1222] = 8'hBC; frame2.valid[1222] = 1'b1; frame2.error[1222] = 1'b0;frame2.data[1223] = 8'hBD; frame2.valid[1223] = 1'b1; frame2.error[1223] = 1'b0;frame2.data[1224] = 8'hBE; frame2.valid[1224] = 1'b1; frame2.error[1224] = 1'b0;frame2.data[1225] = 8'hBF; frame2.valid[1225] = 1'b1; frame2.error[1225] = 1'b0;frame2.data[1226] = 8'hC0; frame2.valid[1226] = 1'b1; frame2.error[1226] = 1'b0;frame2.data[1227] = 8'hC1; frame2.valid[1227] = 1'b1; frame2.error[1227] = 1'b0;frame2.data[1228] = 8'hC2; frame2.valid[1228] = 1'b1; frame2.error[1228] = 1'b0;frame2.data[1229] = 8'hC3; frame2.valid[1229] = 1'b1; frame2.error[1229] = 1'b0;
        frame2.data[1230] = 8'hC4; frame2.valid[1230] = 1'b1; frame2.error[1230] = 1'b0;frame2.data[1231] = 8'hC5; frame2.valid[1231] = 1'b1; frame2.error[1231] = 1'b0;frame2.data[1232] = 8'hC6; frame2.valid[1232] = 1'b1; frame2.error[1232] = 1'b0;frame2.data[1233] = 8'hC7; frame2.valid[1233] = 1'b1; frame2.error[1233] = 1'b0;frame2.data[1234] = 8'hC8; frame2.valid[1234] = 1'b1; frame2.error[1234] = 1'b0;frame2.data[1235] = 8'hC9; frame2.valid[1235] = 1'b1; frame2.error[1235] = 1'b0;frame2.data[1236] = 8'hCA; frame2.valid[1236] = 1'b1; frame2.error[1236] = 1'b0;frame2.data[1237] = 8'hCB; frame2.valid[1237] = 1'b1; frame2.error[1237] = 1'b0;frame2.data[1238] = 8'hCC; frame2.valid[1238] = 1'b1; frame2.error[1238] = 1'b0;frame2.data[1239] = 8'hCD; frame2.valid[1239] = 1'b1; frame2.error[1239] = 1'b0;frame2.data[1240] = 8'hCE; frame2.valid[1240] = 1'b1; frame2.error[1240] = 1'b0;frame2.data[1241] = 8'hCF; frame2.valid[1241] = 1'b1; frame2.error[1241] = 1'b0;frame2.data[1242] = 8'hD0; frame2.valid[1242] = 1'b1; frame2.error[1242] = 1'b0;frame2.data[1243] = 8'hD1; frame2.valid[1243] = 1'b1; frame2.error[1243] = 1'b0;frame2.data[1244] = 8'hD2; frame2.valid[1244] = 1'b1; frame2.error[1244] = 1'b0;frame2.data[1245] = 8'hD3; frame2.valid[1245] = 1'b1; frame2.error[1245] = 1'b0;
        frame2.data[1246] = 8'hD4; frame2.valid[1246] = 1'b1; frame2.error[1246] = 1'b0;frame2.data[1247] = 8'hD5; frame2.valid[1247] = 1'b1; frame2.error[1247] = 1'b0;frame2.data[1248] = 8'hD6; frame2.valid[1248] = 1'b1; frame2.error[1248] = 1'b0;frame2.data[1249] = 8'hD7; frame2.valid[1249] = 1'b1; frame2.error[1249] = 1'b0;frame2.data[1250] = 8'hD8; frame2.valid[1250] = 1'b1; frame2.error[1250] = 1'b0;frame2.data[1251] = 8'hD9; frame2.valid[1251] = 1'b1; frame2.error[1251] = 1'b0;frame2.data[1252] = 8'hDA; frame2.valid[1252] = 1'b1; frame2.error[1252] = 1'b0;frame2.data[1253] = 8'hDB; frame2.valid[1253] = 1'b1; frame2.error[1253] = 1'b0;frame2.data[1254] = 8'hDC; frame2.valid[1254] = 1'b1; frame2.error[1254] = 1'b0;frame2.data[1255] = 8'hDD; frame2.valid[1255] = 1'b1; frame2.error[1255] = 1'b0;frame2.data[1256] = 8'hDE; frame2.valid[1256] = 1'b1; frame2.error[1256] = 1'b0;frame2.data[1257] = 8'hDF; frame2.valid[1257] = 1'b1; frame2.error[1257] = 1'b0;frame2.data[1258] = 8'hE0; frame2.valid[1258] = 1'b1; frame2.error[1258] = 1'b0;frame2.data[1259] = 8'hE1; frame2.valid[1259] = 1'b1; frame2.error[1259] = 1'b0;frame2.data[1260] = 8'hE2; frame2.valid[1260] = 1'b1; frame2.error[1260] = 1'b0;frame2.data[1261] = 8'hE3; frame2.valid[1261] = 1'b1; frame2.error[1261] = 1'b0;
        frame2.data[1262] = 8'hE4; frame2.valid[1262] = 1'b1; frame2.error[1262] = 1'b0;frame2.data[1263] = 8'hE5; frame2.valid[1263] = 1'b1; frame2.error[1263] = 1'b0;frame2.data[1264] = 8'hE6; frame2.valid[1264] = 1'b1; frame2.error[1264] = 1'b0;frame2.data[1265] = 8'hE7; frame2.valid[1265] = 1'b1; frame2.error[1265] = 1'b0;frame2.data[1266] = 8'hE8; frame2.valid[1266] = 1'b1; frame2.error[1266] = 1'b0;frame2.data[1267] = 8'hE9; frame2.valid[1267] = 1'b1; frame2.error[1267] = 1'b0;frame2.data[1268] = 8'hEA; frame2.valid[1268] = 1'b1; frame2.error[1268] = 1'b0;frame2.data[1269] = 8'hEB; frame2.valid[1269] = 1'b1; frame2.error[1269] = 1'b0;frame2.data[1270] = 8'hEC; frame2.valid[1270] = 1'b1; frame2.error[1270] = 1'b0;frame2.data[1271] = 8'hED; frame2.valid[1271] = 1'b1; frame2.error[1271] = 1'b0;frame2.data[1272] = 8'hEE; frame2.valid[1272] = 1'b1; frame2.error[1272] = 1'b0;frame2.data[1273] = 8'hEF; frame2.valid[1273] = 1'b1; frame2.error[1273] = 1'b0;frame2.data[1274] = 8'hF0; frame2.valid[1274] = 1'b1; frame2.error[1274] = 1'b0;frame2.data[1275] = 8'hF1; frame2.valid[1275] = 1'b1; frame2.error[1275] = 1'b0;frame2.data[1276] = 8'hF2; frame2.valid[1276] = 1'b1; frame2.error[1276] = 1'b0;frame2.data[1277] = 8'hF3; frame2.valid[1277] = 1'b1; frame2.error[1277] = 1'b0;
        frame2.data[1278] = 8'hF4; frame2.valid[1278] = 1'b1; frame2.error[1278] = 1'b0;frame2.data[1279] = 8'hF5; frame2.valid[1279] = 1'b1; frame2.error[1279] = 1'b0;frame2.data[1280] = 8'hF6; frame2.valid[1280] = 1'b1; frame2.error[1280] = 1'b0;frame2.data[1281] = 8'hF7; frame2.valid[1281] = 1'b1; frame2.error[1281] = 1'b0;frame2.data[1282] = 8'hF8; frame2.valid[1282] = 1'b1; frame2.error[1282] = 1'b0;frame2.data[1283] = 8'hF9; frame2.valid[1283] = 1'b1; frame2.error[1283] = 1'b0;frame2.data[1284] = 8'hFA; frame2.valid[1284] = 1'b1; frame2.error[1284] = 1'b0;frame2.data[1285] = 8'hFB; frame2.valid[1285] = 1'b1; frame2.error[1285] = 1'b0;frame2.data[1286] = 8'hFC; frame2.valid[1286] = 1'b1; frame2.error[1286] = 1'b0;frame2.data[1287] = 8'hFD; frame2.valid[1287] = 1'b1; frame2.error[1287] = 1'b0;frame2.data[1288] = 8'hFE; frame2.valid[1288] = 1'b1; frame2.error[1288] = 1'b0;frame2.data[1289] = 8'h00; frame2.valid[1289] = 1'b1; frame2.error[1289] = 1'b0;frame2.data[1290] = 8'h01; frame2.valid[1290] = 1'b1; frame2.error[1290] = 1'b0;frame2.data[1291] = 8'h02; frame2.valid[1291] = 1'b1; frame2.error[1291] = 1'b0;frame2.data[1292] = 8'h03; frame2.valid[1292] = 1'b1; frame2.error[1292] = 1'b0;frame2.data[1293] = 8'h04; frame2.valid[1293] = 1'b1; frame2.error[1293] = 1'b0;
        frame2.data[1294] = 8'h05; frame2.valid[1294] = 1'b1; frame2.error[1294] = 1'b0;frame2.data[1295] = 8'h06; frame2.valid[1295] = 1'b1; frame2.error[1295] = 1'b0;frame2.data[1296] = 8'h07; frame2.valid[1296] = 1'b1; frame2.error[1296] = 1'b0;frame2.data[1297] = 8'h08; frame2.valid[1297] = 1'b1; frame2.error[1297] = 1'b0;frame2.data[1298] = 8'h09; frame2.valid[1298] = 1'b1; frame2.error[1298] = 1'b0;frame2.data[1299] = 8'h0A; frame2.valid[1299] = 1'b1; frame2.error[1299] = 1'b0;frame2.data[1300] = 8'h0B; frame2.valid[1300] = 1'b1; frame2.error[1300] = 1'b0;frame2.data[1301] = 8'h0C; frame2.valid[1301] = 1'b1; frame2.error[1301] = 1'b0;frame2.data[1302] = 8'h0D; frame2.valid[1302] = 1'b1; frame2.error[1302] = 1'b0;frame2.data[1303] = 8'h0E; frame2.valid[1303] = 1'b1; frame2.error[1303] = 1'b0;frame2.data[1304] = 8'h0F; frame2.valid[1304] = 1'b1; frame2.error[1304] = 1'b0;frame2.data[1305] = 8'h10; frame2.valid[1305] = 1'b1; frame2.error[1305] = 1'b0;frame2.data[1306] = 8'h11; frame2.valid[1306] = 1'b1; frame2.error[1306] = 1'b0;frame2.data[1307] = 8'h12; frame2.valid[1307] = 1'b1; frame2.error[1307] = 1'b0;frame2.data[1308] = 8'h13; frame2.valid[1308] = 1'b1; frame2.error[1308] = 1'b0;frame2.data[1309] = 8'h14; frame2.valid[1309] = 1'b1; frame2.error[1309] = 1'b0;
        frame2.data[1310] = 8'h15; frame2.valid[1310] = 1'b1; frame2.error[1310] = 1'b0;frame2.data[1311] = 8'h16; frame2.valid[1311] = 1'b1; frame2.error[1311] = 1'b0;frame2.data[1312] = 8'h17; frame2.valid[1312] = 1'b1; frame2.error[1312] = 1'b0;frame2.data[1313] = 8'h18; frame2.valid[1313] = 1'b1; frame2.error[1313] = 1'b0;frame2.data[1314] = 8'h19; frame2.valid[1314] = 1'b1; frame2.error[1314] = 1'b0;frame2.data[1315] = 8'h1A; frame2.valid[1315] = 1'b1; frame2.error[1315] = 1'b0;frame2.data[1316] = 8'h1B; frame2.valid[1316] = 1'b1; frame2.error[1316] = 1'b0;frame2.data[1317] = 8'h1C; frame2.valid[1317] = 1'b1; frame2.error[1317] = 1'b0;frame2.data[1318] = 8'h1D; frame2.valid[1318] = 1'b1; frame2.error[1318] = 1'b0;frame2.data[1319] = 8'h1E; frame2.valid[1319] = 1'b1; frame2.error[1319] = 1'b0;frame2.data[1320] = 8'h1F; frame2.valid[1320] = 1'b1; frame2.error[1320] = 1'b0;frame2.data[1321] = 8'h20; frame2.valid[1321] = 1'b1; frame2.error[1321] = 1'b0;frame2.data[1322] = 8'h21; frame2.valid[1322] = 1'b1; frame2.error[1322] = 1'b0;frame2.data[1323] = 8'h22; frame2.valid[1323] = 1'b1; frame2.error[1323] = 1'b0;frame2.data[1324] = 8'h23; frame2.valid[1324] = 1'b1; frame2.error[1324] = 1'b0;frame2.data[1325] = 8'h24; frame2.valid[1325] = 1'b1; frame2.error[1325] = 1'b0;
        frame2.data[1326] = 8'h25; frame2.valid[1326] = 1'b1; frame2.error[1326] = 1'b0;frame2.data[1327] = 8'h26; frame2.valid[1327] = 1'b1; frame2.error[1327] = 1'b0;frame2.data[1328] = 8'h27; frame2.valid[1328] = 1'b1; frame2.error[1328] = 1'b0;frame2.data[1329] = 8'h28; frame2.valid[1329] = 1'b1; frame2.error[1329] = 1'b0;frame2.data[1330] = 8'h29; frame2.valid[1330] = 1'b1; frame2.error[1330] = 1'b0;frame2.data[1331] = 8'h2A; frame2.valid[1331] = 1'b1; frame2.error[1331] = 1'b0;frame2.data[1332] = 8'h2B; frame2.valid[1332] = 1'b1; frame2.error[1332] = 1'b0;frame2.data[1333] = 8'h2C; frame2.valid[1333] = 1'b1; frame2.error[1333] = 1'b0;frame2.data[1334] = 8'h2D; frame2.valid[1334] = 1'b1; frame2.error[1334] = 1'b0;frame2.data[1335] = 8'h2E; frame2.valid[1335] = 1'b1; frame2.error[1335] = 1'b0;frame2.data[1336] = 8'h2F; frame2.valid[1336] = 1'b1; frame2.error[1336] = 1'b0;frame2.data[1337] = 8'h30; frame2.valid[1337] = 1'b1; frame2.error[1337] = 1'b0;frame2.data[1338] = 8'h31; frame2.valid[1338] = 1'b1; frame2.error[1338] = 1'b0;frame2.data[1339] = 8'h32; frame2.valid[1339] = 1'b1; frame2.error[1339] = 1'b0;frame2.data[1340] = 8'h33; frame2.valid[1340] = 1'b1; frame2.error[1340] = 1'b0;frame2.data[1341] = 8'h34; frame2.valid[1341] = 1'b1; frame2.error[1341] = 1'b0;
        frame2.data[1342] = 8'h35; frame2.valid[1342] = 1'b1; frame2.error[1342] = 1'b0;frame2.data[1343] = 8'h36; frame2.valid[1343] = 1'b1; frame2.error[1343] = 1'b0;frame2.data[1344] = 8'h37; frame2.valid[1344] = 1'b1; frame2.error[1344] = 1'b0;frame2.data[1345] = 8'h38; frame2.valid[1345] = 1'b1; frame2.error[1345] = 1'b0;frame2.data[1346] = 8'h39; frame2.valid[1346] = 1'b1; frame2.error[1346] = 1'b0;frame2.data[1347] = 8'h3A; frame2.valid[1347] = 1'b1; frame2.error[1347] = 1'b0;frame2.data[1348] = 8'h3B; frame2.valid[1348] = 1'b1; frame2.error[1348] = 1'b0;frame2.data[1349] = 8'h3C; frame2.valid[1349] = 1'b1; frame2.error[1349] = 1'b0;frame2.data[1350] = 8'h3D; frame2.valid[1350] = 1'b1; frame2.error[1350] = 1'b0;frame2.data[1351] = 8'h3E; frame2.valid[1351] = 1'b1; frame2.error[1351] = 1'b0;frame2.data[1352] = 8'h3F; frame2.valid[1352] = 1'b1; frame2.error[1352] = 1'b0;frame2.data[1353] = 8'h40; frame2.valid[1353] = 1'b1; frame2.error[1353] = 1'b0;frame2.data[1354] = 8'h41; frame2.valid[1354] = 1'b1; frame2.error[1354] = 1'b0;frame2.data[1355] = 8'h42; frame2.valid[1355] = 1'b1; frame2.error[1355] = 1'b0;frame2.data[1356] = 8'h43; frame2.valid[1356] = 1'b1; frame2.error[1356] = 1'b0;frame2.data[1357] = 8'h44; frame2.valid[1357] = 1'b1; frame2.error[1357] = 1'b0;
        frame2.data[1358] = 8'h45; frame2.valid[1358] = 1'b1; frame2.error[1358] = 1'b0;frame2.data[1359] = 8'h46; frame2.valid[1359] = 1'b1; frame2.error[1359] = 1'b0;frame2.data[1360] = 8'h47; frame2.valid[1360] = 1'b1; frame2.error[1360] = 1'b0;frame2.data[1361] = 8'h48; frame2.valid[1361] = 1'b1; frame2.error[1361] = 1'b0;frame2.data[1362] = 8'h49; frame2.valid[1362] = 1'b1; frame2.error[1362] = 1'b0;frame2.data[1363] = 8'h4A; frame2.valid[1363] = 1'b1; frame2.error[1363] = 1'b0;frame2.data[1364] = 8'h4B; frame2.valid[1364] = 1'b1; frame2.error[1364] = 1'b0;frame2.data[1365] = 8'h4C; frame2.valid[1365] = 1'b1; frame2.error[1365] = 1'b0;frame2.data[1366] = 8'h4D; frame2.valid[1366] = 1'b1; frame2.error[1366] = 1'b0;frame2.data[1367] = 8'h4E; frame2.valid[1367] = 1'b1; frame2.error[1367] = 1'b0;frame2.data[1368] = 8'h4F; frame2.valid[1368] = 1'b1; frame2.error[1368] = 1'b0;frame2.data[1369] = 8'h50; frame2.valid[1369] = 1'b1; frame2.error[1369] = 1'b0;frame2.data[1370] = 8'h51; frame2.valid[1370] = 1'b1; frame2.error[1370] = 1'b0;frame2.data[1371] = 8'h52; frame2.valid[1371] = 1'b1; frame2.error[1371] = 1'b0;frame2.data[1372] = 8'h53; frame2.valid[1372] = 1'b1; frame2.error[1372] = 1'b0;frame2.data[1373] = 8'h54; frame2.valid[1373] = 1'b1; frame2.error[1373] = 1'b0;
        frame2.data[1374] = 8'h55; frame2.valid[1374] = 1'b1; frame2.error[1374] = 1'b0;frame2.data[1375] = 8'h56; frame2.valid[1375] = 1'b1; frame2.error[1375] = 1'b0;frame2.data[1376] = 8'h57; frame2.valid[1376] = 1'b1; frame2.error[1376] = 1'b0;frame2.data[1377] = 8'h58; frame2.valid[1377] = 1'b1; frame2.error[1377] = 1'b0;frame2.data[1378] = 8'h59; frame2.valid[1378] = 1'b1; frame2.error[1378] = 1'b0;frame2.data[1379] = 8'h5A; frame2.valid[1379] = 1'b1; frame2.error[1379] = 1'b0;frame2.data[1380] = 8'h5B; frame2.valid[1380] = 1'b1; frame2.error[1380] = 1'b0;frame2.data[1381] = 8'h5C; frame2.valid[1381] = 1'b1; frame2.error[1381] = 1'b0;frame2.data[1382] = 8'h5D; frame2.valid[1382] = 1'b1; frame2.error[1382] = 1'b0;frame2.data[1383] = 8'h5E; frame2.valid[1383] = 1'b1; frame2.error[1383] = 1'b0;frame2.data[1384] = 8'h5F; frame2.valid[1384] = 1'b1; frame2.error[1384] = 1'b0;frame2.data[1385] = 8'h60; frame2.valid[1385] = 1'b1; frame2.error[1385] = 1'b0;frame2.data[1386] = 8'h61; frame2.valid[1386] = 1'b1; frame2.error[1386] = 1'b0;frame2.data[1387] = 8'h62; frame2.valid[1387] = 1'b1; frame2.error[1387] = 1'b0;frame2.data[1388] = 8'h63; frame2.valid[1388] = 1'b1; frame2.error[1388] = 1'b0;frame2.data[1389] = 8'h64; frame2.valid[1389] = 1'b1; frame2.error[1389] = 1'b0;
        frame2.data[1390] = 8'h65; frame2.valid[1390] = 1'b1; frame2.error[1390] = 1'b0;frame2.data[1391] = 8'h66; frame2.valid[1391] = 1'b1; frame2.error[1391] = 1'b0;frame2.data[1392] = 8'h67; frame2.valid[1392] = 1'b1; frame2.error[1392] = 1'b0;frame2.data[1393] = 8'h68; frame2.valid[1393] = 1'b1; frame2.error[1393] = 1'b0;frame2.data[1394] = 8'h69; frame2.valid[1394] = 1'b1; frame2.error[1394] = 1'b0;frame2.data[1395] = 8'h6A; frame2.valid[1395] = 1'b1; frame2.error[1395] = 1'b0;frame2.data[1396] = 8'h6B; frame2.valid[1396] = 1'b1; frame2.error[1396] = 1'b0;frame2.data[1397] = 8'h6C; frame2.valid[1397] = 1'b1; frame2.error[1397] = 1'b0;frame2.data[1398] = 8'h6D; frame2.valid[1398] = 1'b1; frame2.error[1398] = 1'b0;frame2.data[1399] = 8'h6E; frame2.valid[1399] = 1'b1; frame2.error[1399] = 1'b0;frame2.data[1400] = 8'h6F; frame2.valid[1400] = 1'b1; frame2.error[1400] = 1'b0;frame2.data[1401] = 8'h70; frame2.valid[1401] = 1'b1; frame2.error[1401] = 1'b0;frame2.data[1402] = 8'h71; frame2.valid[1402] = 1'b1; frame2.error[1402] = 1'b0;frame2.data[1403] = 8'h72; frame2.valid[1403] = 1'b1; frame2.error[1403] = 1'b0;frame2.data[1404] = 8'h73; frame2.valid[1404] = 1'b1; frame2.error[1404] = 1'b0;frame2.data[1405] = 8'h74; frame2.valid[1405] = 1'b1; frame2.error[1405] = 1'b0;
        frame2.data[1406] = 8'h75; frame2.valid[1406] = 1'b1; frame2.error[1406] = 1'b0;frame2.data[1407] = 8'h76; frame2.valid[1407] = 1'b1; frame2.error[1407] = 1'b0;frame2.data[1408] = 8'h77; frame2.valid[1408] = 1'b1; frame2.error[1408] = 1'b0;frame2.data[1409] = 8'h78; frame2.valid[1409] = 1'b1; frame2.error[1409] = 1'b0;frame2.data[1410] = 8'h79; frame2.valid[1410] = 1'b1; frame2.error[1410] = 1'b0;frame2.data[1411] = 8'h7A; frame2.valid[1411] = 1'b1; frame2.error[1411] = 1'b0;frame2.data[1412] = 8'h7B; frame2.valid[1412] = 1'b1; frame2.error[1412] = 1'b0;frame2.data[1413] = 8'h7C; frame2.valid[1413] = 1'b1; frame2.error[1413] = 1'b0;frame2.data[1414] = 8'h7D; frame2.valid[1414] = 1'b1; frame2.error[1414] = 1'b0;frame2.data[1415] = 8'h7E; frame2.valid[1415] = 1'b1; frame2.error[1415] = 1'b0;frame2.data[1416] = 8'h7F; frame2.valid[1416] = 1'b1; frame2.error[1416] = 1'b0;frame2.data[1417] = 8'h80; frame2.valid[1417] = 1'b1; frame2.error[1417] = 1'b0;frame2.data[1418] = 8'h81; frame2.valid[1418] = 1'b1; frame2.error[1418] = 1'b0;frame2.data[1419] = 8'h82; frame2.valid[1419] = 1'b1; frame2.error[1419] = 1'b0;frame2.data[1420] = 8'h83; frame2.valid[1420] = 1'b1; frame2.error[1420] = 1'b0;frame2.data[1421] = 8'h84; frame2.valid[1421] = 1'b1; frame2.error[1421] = 1'b0;
        frame2.data[1422] = 8'h85; frame2.valid[1422] = 1'b1; frame2.error[1422] = 1'b0;frame2.data[1423] = 8'h86; frame2.valid[1423] = 1'b1; frame2.error[1423] = 1'b0;frame2.data[1424] = 8'h87; frame2.valid[1424] = 1'b1; frame2.error[1424] = 1'b0;frame2.data[1425] = 8'h88; frame2.valid[1425] = 1'b1; frame2.error[1425] = 1'b0;frame2.data[1426] = 8'h89; frame2.valid[1426] = 1'b1; frame2.error[1426] = 1'b0;frame2.data[1427] = 8'h8A; frame2.valid[1427] = 1'b1; frame2.error[1427] = 1'b0;frame2.data[1428] = 8'h8B; frame2.valid[1428] = 1'b1; frame2.error[1428] = 1'b0;frame2.data[1429] = 8'h8C; frame2.valid[1429] = 1'b1; frame2.error[1429] = 1'b0;frame2.data[1430] = 8'h8D; frame2.valid[1430] = 1'b1; frame2.error[1430] = 1'b0;frame2.data[1431] = 8'h8E; frame2.valid[1431] = 1'b1; frame2.error[1431] = 1'b0;frame2.data[1432] = 8'h8F; frame2.valid[1432] = 1'b1; frame2.error[1432] = 1'b0;frame2.data[1433] = 8'h90; frame2.valid[1433] = 1'b1; frame2.error[1433] = 1'b0;frame2.data[1434] = 8'h91; frame2.valid[1434] = 1'b1; frame2.error[1434] = 1'b0;frame2.data[1435] = 8'h92; frame2.valid[1435] = 1'b1; frame2.error[1435] = 1'b0;frame2.data[1436] = 8'h93; frame2.valid[1436] = 1'b1; frame2.error[1436] = 1'b0;frame2.data[1437] = 8'h94; frame2.valid[1437] = 1'b1; frame2.error[1437] = 1'b0;
        frame2.data[1438] = 8'h95; frame2.valid[1438] = 1'b1; frame2.error[1438] = 1'b0;frame2.data[1439] = 8'h96; frame2.valid[1439] = 1'b1; frame2.error[1439] = 1'b0;frame2.data[1440] = 8'h97; frame2.valid[1440] = 1'b1; frame2.error[1440] = 1'b0;frame2.data[1441] = 8'h98; frame2.valid[1441] = 1'b1; frame2.error[1441] = 1'b0;frame2.data[1442] = 8'h99; frame2.valid[1442] = 1'b1; frame2.error[1442] = 1'b0;frame2.data[1443] = 8'h9A; frame2.valid[1443] = 1'b1; frame2.error[1443] = 1'b0;frame2.data[1444] = 8'h9B; frame2.valid[1444] = 1'b1; frame2.error[1444] = 1'b0;frame2.data[1445] = 8'h9C; frame2.valid[1445] = 1'b1; frame2.error[1445] = 1'b0;frame2.data[1446] = 8'h9D; frame2.valid[1446] = 1'b1; frame2.error[1446] = 1'b0;frame2.data[1447] = 8'h9E; frame2.valid[1447] = 1'b1; frame2.error[1447] = 1'b0;frame2.data[1448] = 8'h9F; frame2.valid[1448] = 1'b1; frame2.error[1448] = 1'b0;frame2.data[1449] = 8'hA0; frame2.valid[1449] = 1'b1; frame2.error[1449] = 1'b0;frame2.data[1450] = 8'hA1; frame2.valid[1450] = 1'b1; frame2.error[1450] = 1'b0;frame2.data[1451] = 8'hA2; frame2.valid[1451] = 1'b1; frame2.error[1451] = 1'b0;frame2.data[1452] = 8'hA3; frame2.valid[1452] = 1'b1; frame2.error[1452] = 1'b0;frame2.data[1453] = 8'hA4; frame2.valid[1453] = 1'b1; frame2.error[1453] = 1'b0;
        frame2.data[1454] = 8'hA5; frame2.valid[1454] = 1'b1; frame2.error[1454] = 1'b0;frame2.data[1455] = 8'hA6; frame2.valid[1455] = 1'b1; frame2.error[1455] = 1'b0;frame2.data[1456] = 8'hA7; frame2.valid[1456] = 1'b1; frame2.error[1456] = 1'b0;frame2.data[1457] = 8'hA8; frame2.valid[1457] = 1'b1; frame2.error[1457] = 1'b0;frame2.data[1458] = 8'hA9; frame2.valid[1458] = 1'b1; frame2.error[1458] = 1'b0;frame2.data[1459] = 8'hAA; frame2.valid[1459] = 1'b1; frame2.error[1459] = 1'b0;frame2.data[1460] = 8'hAB; frame2.valid[1460] = 1'b1; frame2.error[1460] = 1'b0;frame2.data[1461] = 8'hAC; frame2.valid[1461] = 1'b1; frame2.error[1461] = 1'b0;frame2.data[1462] = 8'hAD; frame2.valid[1462] = 1'b1; frame2.error[1462] = 1'b0;frame2.data[1463] = 8'hAE; frame2.valid[1463] = 1'b1; frame2.error[1463] = 1'b0;frame2.data[1464] = 8'hAF; frame2.valid[1464] = 1'b1; frame2.error[1464] = 1'b0;frame2.data[1465] = 8'hB0; frame2.valid[1465] = 1'b1; frame2.error[1465] = 1'b0;frame2.data[1466] = 8'hB1; frame2.valid[1466] = 1'b1; frame2.error[1466] = 1'b0;frame2.data[1467] = 8'hB2; frame2.valid[1467] = 1'b1; frame2.error[1467] = 1'b0;frame2.data[1468] = 8'hB3; frame2.valid[1468] = 1'b1; frame2.error[1468] = 1'b0;frame2.data[1469] = 8'hB4; frame2.valid[1469] = 1'b1; frame2.error[1469] = 1'b0;
        frame2.data[1470] = 8'hB5; frame2.valid[1470] = 1'b1; frame2.error[1470] = 1'b0;frame2.data[1471] = 8'hB6; frame2.valid[1471] = 1'b1; frame2.error[1471] = 1'b0;frame2.data[1472] = 8'hB7; frame2.valid[1472] = 1'b1; frame2.error[1472] = 1'b0;frame2.data[1473] = 8'hB8; frame2.valid[1473] = 1'b1; frame2.error[1473] = 1'b0;frame2.data[1474] = 8'hB9; frame2.valid[1474] = 1'b1; frame2.error[1474] = 1'b0;frame2.data[1475] = 8'hBA; frame2.valid[1475] = 1'b1; frame2.error[1475] = 1'b0;frame2.data[1476] = 8'hBB; frame2.valid[1476] = 1'b1; frame2.error[1476] = 1'b0;frame2.data[1477] = 8'hBC; frame2.valid[1477] = 1'b1; frame2.error[1477] = 1'b0;frame2.data[1478] = 8'hBD; frame2.valid[1478] = 1'b1; frame2.error[1478] = 1'b0;frame2.data[1479] = 8'hBE; frame2.valid[1479] = 1'b1; frame2.error[1479] = 1'b0;frame2.data[1480] = 8'hBF; frame2.valid[1480] = 1'b1; frame2.error[1480] = 1'b0;frame2.data[1481] = 8'hC0; frame2.valid[1481] = 1'b1; frame2.error[1481] = 1'b0;frame2.data[1482] = 8'hC1; frame2.valid[1482] = 1'b1; frame2.error[1482] = 1'b0;frame2.data[1483] = 8'hC2; frame2.valid[1483] = 1'b1; frame2.error[1483] = 1'b0;frame2.data[1484] = 8'hC3; frame2.valid[1484] = 1'b1; frame2.error[1484] = 1'b0;frame2.data[1485] = 8'hC4; frame2.valid[1485] = 1'b1; frame2.error[1485] = 1'b0;
        frame2.data[1486] = 8'hC5; frame2.valid[1486] = 1'b1; frame2.error[1486] = 1'b0;frame2.data[1487] = 8'hC6; frame2.valid[1487] = 1'b1; frame2.error[1487] = 1'b0;frame2.data[1488] = 8'hC7; frame2.valid[1488] = 1'b1; frame2.error[1488] = 1'b0;frame2.data[1489] = 8'hC8; frame2.valid[1489] = 1'b1; frame2.error[1489] = 1'b0;frame2.data[1490] = 8'hC9; frame2.valid[1490] = 1'b1; frame2.error[1490] = 1'b0;frame2.data[1491] = 8'hCA; frame2.valid[1491] = 1'b1; frame2.error[1491] = 1'b0;frame2.data[1492] = 8'hCB; frame2.valid[1492] = 1'b1; frame2.error[1492] = 1'b0;frame2.data[1493] = 8'hCC; frame2.valid[1493] = 1'b1; frame2.error[1493] = 1'b0;frame2.data[1494] = 8'hCD; frame2.valid[1494] = 1'b1; frame2.error[1494] = 1'b0;frame2.data[1495] = 8'hCE; frame2.valid[1495] = 1'b1; frame2.error[1495] = 1'b0;frame2.data[1496] = 8'hCF; frame2.valid[1496] = 1'b1; frame2.error[1496] = 1'b0;frame2.data[1497] = 8'hD0; frame2.valid[1497] = 1'b1; frame2.error[1497] = 1'b0;frame2.data[1498] = 8'hD1; frame2.valid[1498] = 1'b1; frame2.error[1498] = 1'b0;frame2.data[1499] = 8'hD2; frame2.valid[1499] = 1'b1; frame2.error[1499] = 1'b0;frame2.data[1500] = 8'hD3; frame2.valid[1500] = 1'b1; frame2.error[1500] = 1'b0;frame2.data[1501] = 8'hD4; frame2.valid[1501] = 1'b1; frame2.error[1501] = 1'b0;
        frame2.data[1502] = 8'hD5; frame2.valid[1502] = 1'b1; frame2.error[1502] = 1'b0;frame2.data[1503] = 8'hD6; frame2.valid[1503] = 1'b1; frame2.error[1503] = 1'b0;frame2.data[1504] = 8'hD7; frame2.valid[1504] = 1'b1; frame2.error[1504] = 1'b0;frame2.data[1505] = 8'hD8; frame2.valid[1505] = 1'b1; frame2.error[1505] = 1'b0;frame2.data[1506] = 8'hD9; frame2.valid[1506] = 1'b1; frame2.error[1506] = 1'b0;frame2.data[1507] = 8'hDA; frame2.valid[1507] = 1'b1; frame2.error[1507] = 1'b0;frame2.data[1508] = 8'hDB; frame2.valid[1508] = 1'b1; frame2.error[1508] = 1'b0;frame2.data[1509] = 8'hDC; frame2.valid[1509] = 1'b1; frame2.error[1509] = 1'b0;frame2.data[1510] = 8'hDD; frame2.valid[1510] = 1'b1; frame2.error[1510] = 1'b0;frame2.data[1511] = 8'hDE; frame2.valid[1511] = 1'b1; frame2.error[1511] = 1'b0;frame2.data[1512] = 8'hDF; frame2.valid[1512] = 1'b1; frame2.error[1512] = 1'b0;frame2.data[1513] = 8'hE0; frame2.valid[1513] = 1'b1; frame2.error[1513] = 1'b0;


        frame2.data[1514] = 8'h00;  frame2.valid[1514] = 1'b0;  frame2.error[1514] = 1'b0;
        frame2.data[1515] = 8'h00;  frame2.valid[1515] = 1'b0;  frame2.error[1515] = 1'b0;

        // No error in this frame
        frame2.bad_frame  = 1'b0;

        //-----------
        // Frame 3
        //-----------
        frame3.data[0]  = 8'h00;  frame3.valid[0]  = 1'b1;  frame3.error[0]  = 1'b0; // Destination Address (03)
        frame3.data[1]  = 8'h00;  frame3.valid[1]  = 1'b1;  frame3.error[1]  = 1'b0;
        frame3.data[2]  = 8'h00;  frame3.valid[2]  = 1'b1;  frame3.error[2]  = 1'b0;
        frame3.data[3]  = 8'h00;  frame3.valid[3]  = 1'b1;  frame3.error[3]  = 1'b0;
        frame3.data[4]  = 8'h00;  frame3.valid[4]  = 1'b1;  frame3.error[4]  = 1'b0;
        frame3.data[5]  = 8'h03;  frame3.valid[5]  = 1'b1;  frame3.error[5]  = 1'b0;
        frame3.data[6]  = 8'h00;  frame3.valid[6]  = 1'b1;  frame3.error[6]  = 1'b0; // Source Address  (04)
        frame3.data[7]  = 8'h00;  frame3.valid[7]  = 1'b1;  frame3.error[7]  = 1'b0;
        frame3.data[8]  = 8'h00;  frame3.valid[8]  = 1'b1;  frame3.error[8]  = 1'b0;
        frame3.data[9]  = 8'h00;  frame3.valid[9]  = 1'b1;  frame3.error[9]  = 1'b0;
        frame3.data[10] = 8'h00;  frame3.valid[10] = 1'b1;  frame3.error[10] = 1'b0;
        frame3.data[11] = 8'h04;  frame3.valid[11] = 1'b1;  frame3.error[11] = 1'b0;
        frame3.data[12] = 8'h05;  frame3.valid[12] = 1'b1;  frame3.error[12] = 1'b0;
        frame3.data[13] = 8'hDC;  frame3.valid[13] = 1'b1;  frame3.error[13] = 1'b0; // Length/Type = Length = 1500

        frame3.data[  14] = 8'h00; frame3.valid[  14] = 1'b1; frame3.error[  14] = 1'b0;frame3.data[  15] = 8'h01; frame3.valid[  15] = 1'b1; frame3.error[  15] = 1'b0;frame3.data[  16] = 8'h02; frame3.valid[  16] = 1'b1; frame3.error[  16] = 1'b0;frame3.data[  17] = 8'h03; frame3.valid[  17] = 1'b1; frame3.error[  17] = 1'b0;frame3.data[  18] = 8'h04; frame3.valid[  18] = 1'b1; frame3.error[  18] = 1'b0;frame3.data[  19] = 8'h05; frame3.valid[  19] = 1'b1; frame3.error[  19] = 1'b0;frame3.data[  20] = 8'h06; frame3.valid[  20] = 1'b1; frame3.error[  20] = 1'b0;frame3.data[  21] = 8'h07; frame3.valid[  21] = 1'b1; frame3.error[  21] = 1'b0;frame3.data[  22] = 8'h08; frame3.valid[  22] = 1'b1; frame3.error[  22] = 1'b0;frame3.data[  23] = 8'h09; frame3.valid[  23] = 1'b1; frame3.error[  23] = 1'b0;frame3.data[  24] = 8'h0A; frame3.valid[  24] = 1'b1; frame3.error[  24] = 1'b0;frame3.data[  25] = 8'h0B; frame3.valid[  25] = 1'b1; frame3.error[  25] = 1'b0;frame3.data[  26] = 8'h0C; frame3.valid[  26] = 1'b1; frame3.error[  26] = 1'b0;frame3.data[  27] = 8'h0D; frame3.valid[  27] = 1'b1; frame3.error[  27] = 1'b0;frame3.data[  28] = 8'h0E; frame3.valid[  28] = 1'b1; frame3.error[  28] = 1'b0;frame3.data[  29] = 8'h0F; frame3.valid[  29] = 1'b1; frame3.error[  29] = 1'b0;
        frame3.data[  30] = 8'h10; frame3.valid[  30] = 1'b1; frame3.error[  30] = 1'b0;frame3.data[  31] = 8'h11; frame3.valid[  31] = 1'b1; frame3.error[  31] = 1'b0;frame3.data[  32] = 8'h12; frame3.valid[  32] = 1'b1; frame3.error[  32] = 1'b0;frame3.data[  33] = 8'h13; frame3.valid[  33] = 1'b1; frame3.error[  33] = 1'b0;frame3.data[  34] = 8'h14; frame3.valid[  34] = 1'b1; frame3.error[  34] = 1'b0;frame3.data[  35] = 8'h15; frame3.valid[  35] = 1'b1; frame3.error[  35] = 1'b0;frame3.data[  36] = 8'h16; frame3.valid[  36] = 1'b1; frame3.error[  36] = 1'b0;frame3.data[  37] = 8'h17; frame3.valid[  37] = 1'b1; frame3.error[  37] = 1'b0;frame3.data[  38] = 8'h18; frame3.valid[  38] = 1'b1; frame3.error[  38] = 1'b0;frame3.data[  39] = 8'h19; frame3.valid[  39] = 1'b1; frame3.error[  39] = 1'b0;frame3.data[  40] = 8'h1A; frame3.valid[  40] = 1'b1; frame3.error[  40] = 1'b0;frame3.data[  41] = 8'h1B; frame3.valid[  41] = 1'b1; frame3.error[  41] = 1'b0;frame3.data[  42] = 8'h1C; frame3.valid[  42] = 1'b1; frame3.error[  42] = 1'b0;frame3.data[  43] = 8'h1D; frame3.valid[  43] = 1'b1; frame3.error[  43] = 1'b0;frame3.data[  44] = 8'h1E; frame3.valid[  44] = 1'b1; frame3.error[  44] = 1'b0;frame3.data[  45] = 8'h1F; frame3.valid[  45] = 1'b1; frame3.error[  45] = 1'b0;
        frame3.data[  46] = 8'h20; frame3.valid[  46] = 1'b1; frame3.error[  46] = 1'b0;frame3.data[  47] = 8'h21; frame3.valid[  47] = 1'b1; frame3.error[  47] = 1'b0;frame3.data[  48] = 8'h22; frame3.valid[  48] = 1'b1; frame3.error[  48] = 1'b0;frame3.data[  49] = 8'h23; frame3.valid[  49] = 1'b1; frame3.error[  49] = 1'b0;frame3.data[  50] = 8'h24; frame3.valid[  50] = 1'b1; frame3.error[  50] = 1'b0;frame3.data[  51] = 8'h25; frame3.valid[  51] = 1'b1; frame3.error[  51] = 1'b0;frame3.data[  52] = 8'h26; frame3.valid[  52] = 1'b1; frame3.error[  52] = 1'b0;frame3.data[  53] = 8'h27; frame3.valid[  53] = 1'b1; frame3.error[  53] = 1'b0;frame3.data[  54] = 8'h28; frame3.valid[  54] = 1'b1; frame3.error[  54] = 1'b0;frame3.data[  55] = 8'h29; frame3.valid[  55] = 1'b1; frame3.error[  55] = 1'b0;frame3.data[  56] = 8'h2A; frame3.valid[  56] = 1'b1; frame3.error[  56] = 1'b0;frame3.data[  57] = 8'h2B; frame3.valid[  57] = 1'b1; frame3.error[  57] = 1'b0;frame3.data[  58] = 8'h2C; frame3.valid[  58] = 1'b1; frame3.error[  58] = 1'b0;frame3.data[  59] = 8'h2D; frame3.valid[  59] = 1'b1; frame3.error[  59] = 1'b0;frame3.data[  60] = 8'h2E; frame3.valid[  60] = 1'b1; frame3.error[  60] = 1'b0;frame3.data[  61] = 8'h2F; frame3.valid[  61] = 1'b1; frame3.error[  61] = 1'b0;
        frame3.data[  62] = 8'h30; frame3.valid[  62] = 1'b1; frame3.error[  62] = 1'b0;frame3.data[  63] = 8'h31; frame3.valid[  63] = 1'b1; frame3.error[  63] = 1'b0;frame3.data[  64] = 8'h32; frame3.valid[  64] = 1'b1; frame3.error[  64] = 1'b0;frame3.data[  65] = 8'h33; frame3.valid[  65] = 1'b1; frame3.error[  65] = 1'b0;frame3.data[  66] = 8'h34; frame3.valid[  66] = 1'b1; frame3.error[  66] = 1'b0;frame3.data[  67] = 8'h35; frame3.valid[  67] = 1'b1; frame3.error[  67] = 1'b0;frame3.data[  68] = 8'h36; frame3.valid[  68] = 1'b1; frame3.error[  68] = 1'b0;frame3.data[  69] = 8'h37; frame3.valid[  69] = 1'b1; frame3.error[  69] = 1'b0;frame3.data[  70] = 8'h38; frame3.valid[  70] = 1'b1; frame3.error[  70] = 1'b0;frame3.data[  71] = 8'h39; frame3.valid[  71] = 1'b1; frame3.error[  71] = 1'b0;frame3.data[  72] = 8'h3A; frame3.valid[  72] = 1'b1; frame3.error[  72] = 1'b0;frame3.data[  73] = 8'h3B; frame3.valid[  73] = 1'b1; frame3.error[  73] = 1'b0;frame3.data[  74] = 8'h3C; frame3.valid[  74] = 1'b1; frame3.error[  74] = 1'b0;frame3.data[  75] = 8'h3D; frame3.valid[  75] = 1'b1; frame3.error[  75] = 1'b0;frame3.data[  76] = 8'h3E; frame3.valid[  76] = 1'b1; frame3.error[  76] = 1'b0;frame3.data[  77] = 8'h3F; frame3.valid[  77] = 1'b1; frame3.error[  77] = 1'b0;
        frame3.data[  78] = 8'h40; frame3.valid[  78] = 1'b1; frame3.error[  78] = 1'b0;frame3.data[  79] = 8'h41; frame3.valid[  79] = 1'b1; frame3.error[  79] = 1'b0;frame3.data[  80] = 8'h42; frame3.valid[  80] = 1'b1; frame3.error[  80] = 1'b0;frame3.data[  81] = 8'h43; frame3.valid[  81] = 1'b1; frame3.error[  81] = 1'b0;frame3.data[  82] = 8'h44; frame3.valid[  82] = 1'b1; frame3.error[  82] = 1'b0;frame3.data[  83] = 8'h45; frame3.valid[  83] = 1'b1; frame3.error[  83] = 1'b0;frame3.data[  84] = 8'h46; frame3.valid[  84] = 1'b1; frame3.error[  84] = 1'b0;frame3.data[  85] = 8'h47; frame3.valid[  85] = 1'b1; frame3.error[  85] = 1'b0;frame3.data[  86] = 8'h48; frame3.valid[  86] = 1'b1; frame3.error[  86] = 1'b0;frame3.data[  87] = 8'h49; frame3.valid[  87] = 1'b1; frame3.error[  87] = 1'b0;frame3.data[  88] = 8'h4A; frame3.valid[  88] = 1'b1; frame3.error[  88] = 1'b0;frame3.data[  89] = 8'h4B; frame3.valid[  89] = 1'b1; frame3.error[  89] = 1'b0;frame3.data[  90] = 8'h4C; frame3.valid[  90] = 1'b1; frame3.error[  90] = 1'b0;frame3.data[  91] = 8'h4D; frame3.valid[  91] = 1'b1; frame3.error[  91] = 1'b0;frame3.data[  92] = 8'h4E; frame3.valid[  92] = 1'b1; frame3.error[  92] = 1'b0;frame3.data[  93] = 8'h4F; frame3.valid[  93] = 1'b1; frame3.error[  93] = 1'b0;
        frame3.data[  94] = 8'h50; frame3.valid[  94] = 1'b1; frame3.error[  94] = 1'b0;frame3.data[  95] = 8'h51; frame3.valid[  95] = 1'b1; frame3.error[  95] = 1'b0;frame3.data[  96] = 8'h52; frame3.valid[  96] = 1'b1; frame3.error[  96] = 1'b0;frame3.data[  97] = 8'h53; frame3.valid[  97] = 1'b1; frame3.error[  97] = 1'b0;frame3.data[  98] = 8'h54; frame3.valid[  98] = 1'b1; frame3.error[  98] = 1'b0;frame3.data[  99] = 8'h55; frame3.valid[  99] = 1'b1; frame3.error[  99] = 1'b0;frame3.data[ 100] = 8'h56; frame3.valid[ 100] = 1'b1; frame3.error[ 100] = 1'b0;frame3.data[ 101] = 8'h57; frame3.valid[ 101] = 1'b1; frame3.error[ 101] = 1'b0;frame3.data[ 102] = 8'h58; frame3.valid[ 102] = 1'b1; frame3.error[ 102] = 1'b0;frame3.data[ 103] = 8'h59; frame3.valid[ 103] = 1'b1; frame3.error[ 103] = 1'b0;frame3.data[ 104] = 8'h5A; frame3.valid[ 104] = 1'b1; frame3.error[ 104] = 1'b0;frame3.data[ 105] = 8'h5B; frame3.valid[ 105] = 1'b1; frame3.error[ 105] = 1'b0;frame3.data[ 106] = 8'h5C; frame3.valid[ 106] = 1'b1; frame3.error[ 106] = 1'b0;frame3.data[ 107] = 8'h5D; frame3.valid[ 107] = 1'b1; frame3.error[ 107] = 1'b0;frame3.data[ 108] = 8'h5E; frame3.valid[ 108] = 1'b1; frame3.error[ 108] = 1'b0;frame3.data[ 109] = 8'h5F; frame3.valid[ 109] = 1'b1; frame3.error[ 109] = 1'b0;
        frame3.data[ 110] = 8'h60; frame3.valid[ 110] = 1'b1; frame3.error[ 110] = 1'b0;frame3.data[ 111] = 8'h61; frame3.valid[ 111] = 1'b1; frame3.error[ 111] = 1'b0;frame3.data[ 112] = 8'h62; frame3.valid[ 112] = 1'b1; frame3.error[ 112] = 1'b0;frame3.data[ 113] = 8'h63; frame3.valid[ 113] = 1'b1; frame3.error[ 113] = 1'b0;frame3.data[ 114] = 8'h64; frame3.valid[ 114] = 1'b1; frame3.error[ 114] = 1'b0;frame3.data[ 115] = 8'h65; frame3.valid[ 115] = 1'b1; frame3.error[ 115] = 1'b0;frame3.data[ 116] = 8'h66; frame3.valid[ 116] = 1'b1; frame3.error[ 116] = 1'b0;frame3.data[ 117] = 8'h67; frame3.valid[ 117] = 1'b1; frame3.error[ 117] = 1'b0;frame3.data[ 118] = 8'h68; frame3.valid[ 118] = 1'b1; frame3.error[ 118] = 1'b0;frame3.data[ 119] = 8'h69; frame3.valid[ 119] = 1'b1; frame3.error[ 119] = 1'b0;frame3.data[ 120] = 8'h6A; frame3.valid[ 120] = 1'b1; frame3.error[ 120] = 1'b0;frame3.data[ 121] = 8'h6B; frame3.valid[ 121] = 1'b1; frame3.error[ 121] = 1'b0;frame3.data[ 122] = 8'h6C; frame3.valid[ 122] = 1'b1; frame3.error[ 122] = 1'b0;frame3.data[ 123] = 8'h6D; frame3.valid[ 123] = 1'b1; frame3.error[ 123] = 1'b0;frame3.data[ 124] = 8'h6E; frame3.valid[ 124] = 1'b1; frame3.error[ 124] = 1'b0;frame3.data[ 125] = 8'h6F; frame3.valid[ 125] = 1'b1; frame3.error[ 125] = 1'b0;
        frame3.data[ 126] = 8'h70; frame3.valid[ 126] = 1'b1; frame3.error[ 126] = 1'b0;frame3.data[ 127] = 8'h71; frame3.valid[ 127] = 1'b1; frame3.error[ 127] = 1'b0;frame3.data[ 128] = 8'h72; frame3.valid[ 128] = 1'b1; frame3.error[ 128] = 1'b0;frame3.data[ 129] = 8'h73; frame3.valid[ 129] = 1'b1; frame3.error[ 129] = 1'b0;frame3.data[ 130] = 8'h74; frame3.valid[ 130] = 1'b1; frame3.error[ 130] = 1'b0;frame3.data[ 131] = 8'h75; frame3.valid[ 131] = 1'b1; frame3.error[ 131] = 1'b0;frame3.data[ 132] = 8'h76; frame3.valid[ 132] = 1'b1; frame3.error[ 132] = 1'b0;frame3.data[ 133] = 8'h77; frame3.valid[ 133] = 1'b1; frame3.error[ 133] = 1'b0;frame3.data[ 134] = 8'h78; frame3.valid[ 134] = 1'b1; frame3.error[ 134] = 1'b0;frame3.data[ 135] = 8'h79; frame3.valid[ 135] = 1'b1; frame3.error[ 135] = 1'b0;frame3.data[ 136] = 8'h7A; frame3.valid[ 136] = 1'b1; frame3.error[ 136] = 1'b0;frame3.data[ 137] = 8'h7B; frame3.valid[ 137] = 1'b1; frame3.error[ 137] = 1'b0;frame3.data[ 138] = 8'h7C; frame3.valid[ 138] = 1'b1; frame3.error[ 138] = 1'b0;frame3.data[ 139] = 8'h7D; frame3.valid[ 139] = 1'b1; frame3.error[ 139] = 1'b0;frame3.data[ 140] = 8'h7E; frame3.valid[ 140] = 1'b1; frame3.error[ 140] = 1'b0;frame3.data[ 141] = 8'h7F; frame3.valid[ 141] = 1'b1; frame3.error[ 141] = 1'b0;
        frame3.data[ 142] = 8'h80; frame3.valid[ 142] = 1'b1; frame3.error[ 142] = 1'b0;frame3.data[ 143] = 8'h81; frame3.valid[ 143] = 1'b1; frame3.error[ 143] = 1'b0;frame3.data[ 144] = 8'h82; frame3.valid[ 144] = 1'b1; frame3.error[ 144] = 1'b0;frame3.data[ 145] = 8'h83; frame3.valid[ 145] = 1'b1; frame3.error[ 145] = 1'b0;frame3.data[ 146] = 8'h84; frame3.valid[ 146] = 1'b1; frame3.error[ 146] = 1'b0;frame3.data[ 147] = 8'h85; frame3.valid[ 147] = 1'b1; frame3.error[ 147] = 1'b0;frame3.data[ 148] = 8'h86; frame3.valid[ 148] = 1'b1; frame3.error[ 148] = 1'b0;frame3.data[ 149] = 8'h87; frame3.valid[ 149] = 1'b1; frame3.error[ 149] = 1'b0;frame3.data[ 150] = 8'h88; frame3.valid[ 150] = 1'b1; frame3.error[ 150] = 1'b0;frame3.data[ 151] = 8'h89; frame3.valid[ 151] = 1'b1; frame3.error[ 151] = 1'b0;frame3.data[ 152] = 8'h8A; frame3.valid[ 152] = 1'b1; frame3.error[ 152] = 1'b0;frame3.data[ 153] = 8'h8B; frame3.valid[ 153] = 1'b1; frame3.error[ 153] = 1'b0;frame3.data[ 154] = 8'h8C; frame3.valid[ 154] = 1'b1; frame3.error[ 154] = 1'b0;frame3.data[ 155] = 8'h8D; frame3.valid[ 155] = 1'b1; frame3.error[ 155] = 1'b0;frame3.data[ 156] = 8'h8E; frame3.valid[ 156] = 1'b1; frame3.error[ 156] = 1'b0;frame3.data[ 157] = 8'h8F; frame3.valid[ 157] = 1'b1; frame3.error[ 157] = 1'b0;
        frame3.data[ 158] = 8'h90; frame3.valid[ 158] = 1'b1; frame3.error[ 158] = 1'b0;frame3.data[ 159] = 8'h91; frame3.valid[ 159] = 1'b1; frame3.error[ 159] = 1'b0;frame3.data[ 160] = 8'h92; frame3.valid[ 160] = 1'b1; frame3.error[ 160] = 1'b0;frame3.data[ 161] = 8'h93; frame3.valid[ 161] = 1'b1; frame3.error[ 161] = 1'b0;frame3.data[ 162] = 8'h94; frame3.valid[ 162] = 1'b1; frame3.error[ 162] = 1'b0;frame3.data[ 163] = 8'h95; frame3.valid[ 163] = 1'b1; frame3.error[ 163] = 1'b0;frame3.data[ 164] = 8'h96; frame3.valid[ 164] = 1'b1; frame3.error[ 164] = 1'b0;frame3.data[ 165] = 8'h97; frame3.valid[ 165] = 1'b1; frame3.error[ 165] = 1'b0;frame3.data[ 166] = 8'h98; frame3.valid[ 166] = 1'b1; frame3.error[ 166] = 1'b0;frame3.data[ 167] = 8'h99; frame3.valid[ 167] = 1'b1; frame3.error[ 167] = 1'b0;frame3.data[ 168] = 8'h9A; frame3.valid[ 168] = 1'b1; frame3.error[ 168] = 1'b0;frame3.data[ 169] = 8'h9B; frame3.valid[ 169] = 1'b1; frame3.error[ 169] = 1'b0;frame3.data[ 170] = 8'h9C; frame3.valid[ 170] = 1'b1; frame3.error[ 170] = 1'b0;frame3.data[ 171] = 8'h9D; frame3.valid[ 171] = 1'b1; frame3.error[ 171] = 1'b0;frame3.data[ 172] = 8'h9E; frame3.valid[ 172] = 1'b1; frame3.error[ 172] = 1'b0;frame3.data[ 173] = 8'h9F; frame3.valid[ 173] = 1'b1; frame3.error[ 173] = 1'b0;
        frame3.data[ 174] = 8'hA0; frame3.valid[ 174] = 1'b1; frame3.error[ 174] = 1'b0;frame3.data[ 175] = 8'hA1; frame3.valid[ 175] = 1'b1; frame3.error[ 175] = 1'b0;frame3.data[ 176] = 8'hA2; frame3.valid[ 176] = 1'b1; frame3.error[ 176] = 1'b0;frame3.data[ 177] = 8'hA3; frame3.valid[ 177] = 1'b1; frame3.error[ 177] = 1'b0;frame3.data[ 178] = 8'hA4; frame3.valid[ 178] = 1'b1; frame3.error[ 178] = 1'b0;frame3.data[ 179] = 8'hA5; frame3.valid[ 179] = 1'b1; frame3.error[ 179] = 1'b0;frame3.data[ 180] = 8'hA6; frame3.valid[ 180] = 1'b1; frame3.error[ 180] = 1'b0;frame3.data[ 181] = 8'hA7; frame3.valid[ 181] = 1'b1; frame3.error[ 181] = 1'b0;frame3.data[ 182] = 8'hA8; frame3.valid[ 182] = 1'b1; frame3.error[ 182] = 1'b0;frame3.data[ 183] = 8'hA9; frame3.valid[ 183] = 1'b1; frame3.error[ 183] = 1'b0;frame3.data[ 184] = 8'hAA; frame3.valid[ 184] = 1'b1; frame3.error[ 184] = 1'b0;frame3.data[ 185] = 8'hAB; frame3.valid[ 185] = 1'b1; frame3.error[ 185] = 1'b0;frame3.data[ 186] = 8'hAC; frame3.valid[ 186] = 1'b1; frame3.error[ 186] = 1'b0;frame3.data[ 187] = 8'hAD; frame3.valid[ 187] = 1'b1; frame3.error[ 187] = 1'b0;frame3.data[ 188] = 8'hAE; frame3.valid[ 188] = 1'b1; frame3.error[ 188] = 1'b0;frame3.data[ 189] = 8'hAF; frame3.valid[ 189] = 1'b1; frame3.error[ 189] = 1'b0;
        frame3.data[ 190] = 8'hB0; frame3.valid[ 190] = 1'b1; frame3.error[ 190] = 1'b0;frame3.data[ 191] = 8'hB1; frame3.valid[ 191] = 1'b1; frame3.error[ 191] = 1'b0;frame3.data[ 192] = 8'hB2; frame3.valid[ 192] = 1'b1; frame3.error[ 192] = 1'b0;frame3.data[ 193] = 8'hB3; frame3.valid[ 193] = 1'b1; frame3.error[ 193] = 1'b0;frame3.data[ 194] = 8'hB4; frame3.valid[ 194] = 1'b1; frame3.error[ 194] = 1'b0;frame3.data[ 195] = 8'hB5; frame3.valid[ 195] = 1'b1; frame3.error[ 195] = 1'b0;frame3.data[ 196] = 8'hB6; frame3.valid[ 196] = 1'b1; frame3.error[ 196] = 1'b0;frame3.data[ 197] = 8'hB7; frame3.valid[ 197] = 1'b1; frame3.error[ 197] = 1'b0;frame3.data[ 198] = 8'hB8; frame3.valid[ 198] = 1'b1; frame3.error[ 198] = 1'b0;frame3.data[ 199] = 8'hB9; frame3.valid[ 199] = 1'b1; frame3.error[ 199] = 1'b0;frame3.data[ 200] = 8'hBA; frame3.valid[ 200] = 1'b1; frame3.error[ 200] = 1'b0;frame3.data[ 201] = 8'hBB; frame3.valid[ 201] = 1'b1; frame3.error[ 201] = 1'b0;frame3.data[ 202] = 8'hBC; frame3.valid[ 202] = 1'b1; frame3.error[ 202] = 1'b0;frame3.data[ 203] = 8'hBD; frame3.valid[ 203] = 1'b1; frame3.error[ 203] = 1'b0;frame3.data[ 204] = 8'hBE; frame3.valid[ 204] = 1'b1; frame3.error[ 204] = 1'b0;frame3.data[ 205] = 8'hBF; frame3.valid[ 205] = 1'b1; frame3.error[ 205] = 1'b0;
        frame3.data[ 206] = 8'hC0; frame3.valid[ 206] = 1'b1; frame3.error[ 206] = 1'b0;frame3.data[ 207] = 8'hC1; frame3.valid[ 207] = 1'b1; frame3.error[ 207] = 1'b0;frame3.data[ 208] = 8'hC2; frame3.valid[ 208] = 1'b1; frame3.error[ 208] = 1'b0;frame3.data[ 209] = 8'hC3; frame3.valid[ 209] = 1'b1; frame3.error[ 209] = 1'b0;frame3.data[ 210] = 8'hC4; frame3.valid[ 210] = 1'b1; frame3.error[ 210] = 1'b0;frame3.data[ 211] = 8'hC5; frame3.valid[ 211] = 1'b1; frame3.error[ 211] = 1'b0;frame3.data[ 212] = 8'hC6; frame3.valid[ 212] = 1'b1; frame3.error[ 212] = 1'b0;frame3.data[ 213] = 8'hC7; frame3.valid[ 213] = 1'b1; frame3.error[ 213] = 1'b0;frame3.data[ 214] = 8'hC8; frame3.valid[ 214] = 1'b1; frame3.error[ 214] = 1'b0;frame3.data[ 215] = 8'hC9; frame3.valid[ 215] = 1'b1; frame3.error[ 215] = 1'b0;frame3.data[ 216] = 8'hCA; frame3.valid[ 216] = 1'b1; frame3.error[ 216] = 1'b0;frame3.data[ 217] = 8'hCB; frame3.valid[ 217] = 1'b1; frame3.error[ 217] = 1'b0;frame3.data[ 218] = 8'hCC; frame3.valid[ 218] = 1'b1; frame3.error[ 218] = 1'b0;frame3.data[ 219] = 8'hCD; frame3.valid[ 219] = 1'b1; frame3.error[ 219] = 1'b0;frame3.data[ 220] = 8'hCE; frame3.valid[ 220] = 1'b1; frame3.error[ 220] = 1'b0;frame3.data[ 221] = 8'hCF; frame3.valid[ 221] = 1'b1; frame3.error[ 221] = 1'b0;
        frame3.data[ 222] = 8'hD0; frame3.valid[ 222] = 1'b1; frame3.error[ 222] = 1'b0;frame3.data[ 223] = 8'hD1; frame3.valid[ 223] = 1'b1; frame3.error[ 223] = 1'b0;frame3.data[ 224] = 8'hD2; frame3.valid[ 224] = 1'b1; frame3.error[ 224] = 1'b0;frame3.data[ 225] = 8'hD3; frame3.valid[ 225] = 1'b1; frame3.error[ 225] = 1'b0;frame3.data[ 226] = 8'hD4; frame3.valid[ 226] = 1'b1; frame3.error[ 226] = 1'b0;frame3.data[ 227] = 8'hD5; frame3.valid[ 227] = 1'b1; frame3.error[ 227] = 1'b0;frame3.data[ 228] = 8'hD6; frame3.valid[ 228] = 1'b1; frame3.error[ 228] = 1'b0;frame3.data[ 229] = 8'hD7; frame3.valid[ 229] = 1'b1; frame3.error[ 229] = 1'b0;frame3.data[ 230] = 8'hD8; frame3.valid[ 230] = 1'b1; frame3.error[ 230] = 1'b0;frame3.data[ 231] = 8'hD9; frame3.valid[ 231] = 1'b1; frame3.error[ 231] = 1'b0;frame3.data[ 232] = 8'hDA; frame3.valid[ 232] = 1'b1; frame3.error[ 232] = 1'b0;frame3.data[ 233] = 8'hDB; frame3.valid[ 233] = 1'b1; frame3.error[ 233] = 1'b0;frame3.data[ 234] = 8'hDC; frame3.valid[ 234] = 1'b1; frame3.error[ 234] = 1'b0;frame3.data[ 235] = 8'hDD; frame3.valid[ 235] = 1'b1; frame3.error[ 235] = 1'b0;frame3.data[ 236] = 8'hDE; frame3.valid[ 236] = 1'b1; frame3.error[ 236] = 1'b0;frame3.data[ 237] = 8'hDF; frame3.valid[ 237] = 1'b1; frame3.error[ 237] = 1'b0;
        frame3.data[ 238] = 8'hE0; frame3.valid[ 238] = 1'b1; frame3.error[ 238] = 1'b0;frame3.data[ 239] = 8'hE1; frame3.valid[ 239] = 1'b1; frame3.error[ 239] = 1'b0;frame3.data[ 240] = 8'hE2; frame3.valid[ 240] = 1'b1; frame3.error[ 240] = 1'b0;frame3.data[ 241] = 8'hE3; frame3.valid[ 241] = 1'b1; frame3.error[ 241] = 1'b0;frame3.data[ 242] = 8'hE4; frame3.valid[ 242] = 1'b1; frame3.error[ 242] = 1'b0;frame3.data[ 243] = 8'hE5; frame3.valid[ 243] = 1'b1; frame3.error[ 243] = 1'b0;frame3.data[ 244] = 8'hE6; frame3.valid[ 244] = 1'b1; frame3.error[ 244] = 1'b0;frame3.data[ 245] = 8'hE7; frame3.valid[ 245] = 1'b1; frame3.error[ 245] = 1'b0;frame3.data[ 246] = 8'hE8; frame3.valid[ 246] = 1'b1; frame3.error[ 246] = 1'b0;frame3.data[ 247] = 8'hE9; frame3.valid[ 247] = 1'b1; frame3.error[ 247] = 1'b0;frame3.data[ 248] = 8'hEA; frame3.valid[ 248] = 1'b1; frame3.error[ 248] = 1'b0;frame3.data[ 249] = 8'hEB; frame3.valid[ 249] = 1'b1; frame3.error[ 249] = 1'b0;frame3.data[ 250] = 8'hEC; frame3.valid[ 250] = 1'b1; frame3.error[ 250] = 1'b0;frame3.data[ 251] = 8'hED; frame3.valid[ 251] = 1'b1; frame3.error[ 251] = 1'b0;frame3.data[ 252] = 8'hEE; frame3.valid[ 252] = 1'b1; frame3.error[ 252] = 1'b0;frame3.data[ 253] = 8'hEF; frame3.valid[ 253] = 1'b1; frame3.error[ 253] = 1'b0;
        frame3.data[ 254] = 8'hF0; frame3.valid[ 254] = 1'b1; frame3.error[ 254] = 1'b0;frame3.data[ 255] = 8'hF1; frame3.valid[ 255] = 1'b1; frame3.error[ 255] = 1'b0;frame3.data[ 256] = 8'hF2; frame3.valid[ 256] = 1'b1; frame3.error[ 256] = 1'b0;frame3.data[ 257] = 8'hF3; frame3.valid[ 257] = 1'b1; frame3.error[ 257] = 1'b0;frame3.data[ 258] = 8'hF4; frame3.valid[ 258] = 1'b1; frame3.error[ 258] = 1'b0;frame3.data[ 259] = 8'hF5; frame3.valid[ 259] = 1'b1; frame3.error[ 259] = 1'b0;frame3.data[ 260] = 8'hF6; frame3.valid[ 260] = 1'b1; frame3.error[ 260] = 1'b0;frame3.data[ 261] = 8'hF7; frame3.valid[ 261] = 1'b1; frame3.error[ 261] = 1'b0;frame3.data[ 262] = 8'hF8; frame3.valid[ 262] = 1'b1; frame3.error[ 262] = 1'b0;frame3.data[ 263] = 8'hF9; frame3.valid[ 263] = 1'b1; frame3.error[ 263] = 1'b0;frame3.data[ 264] = 8'hFA; frame3.valid[ 264] = 1'b1; frame3.error[ 264] = 1'b0;frame3.data[ 265] = 8'hFB; frame3.valid[ 265] = 1'b1; frame3.error[ 265] = 1'b0;frame3.data[ 266] = 8'hFC; frame3.valid[ 266] = 1'b1; frame3.error[ 266] = 1'b0;frame3.data[ 267] = 8'hFD; frame3.valid[ 267] = 1'b1; frame3.error[ 267] = 1'b0;frame3.data[ 268] = 8'hFE; frame3.valid[ 268] = 1'b1; frame3.error[ 268] = 1'b0;frame3.data[ 269] = 8'h00; frame3.valid[ 269] = 1'b1; frame3.error[ 269] = 1'b0;
        frame3.data[ 270] = 8'h01; frame3.valid[ 270] = 1'b1; frame3.error[ 270] = 1'b0;frame3.data[ 271] = 8'h02; frame3.valid[ 271] = 1'b1; frame3.error[ 271] = 1'b0;frame3.data[ 272] = 8'h03; frame3.valid[ 272] = 1'b1; frame3.error[ 272] = 1'b0;frame3.data[ 273] = 8'h04; frame3.valid[ 273] = 1'b1; frame3.error[ 273] = 1'b0;frame3.data[ 274] = 8'h05; frame3.valid[ 274] = 1'b1; frame3.error[ 274] = 1'b0;frame3.data[ 275] = 8'h06; frame3.valid[ 275] = 1'b1; frame3.error[ 275] = 1'b0;frame3.data[ 276] = 8'h07; frame3.valid[ 276] = 1'b1; frame3.error[ 276] = 1'b0;frame3.data[ 277] = 8'h08; frame3.valid[ 277] = 1'b1; frame3.error[ 277] = 1'b0;frame3.data[ 278] = 8'h09; frame3.valid[ 278] = 1'b1; frame3.error[ 278] = 1'b0;frame3.data[ 279] = 8'h0A; frame3.valid[ 279] = 1'b1; frame3.error[ 279] = 1'b0;frame3.data[ 280] = 8'h0B; frame3.valid[ 280] = 1'b1; frame3.error[ 280] = 1'b0;frame3.data[ 281] = 8'h0C; frame3.valid[ 281] = 1'b1; frame3.error[ 281] = 1'b0;frame3.data[ 282] = 8'h0D; frame3.valid[ 282] = 1'b1; frame3.error[ 282] = 1'b0;frame3.data[ 283] = 8'h0E; frame3.valid[ 283] = 1'b1; frame3.error[ 283] = 1'b0;frame3.data[ 284] = 8'h0F; frame3.valid[ 284] = 1'b1; frame3.error[ 284] = 1'b0;frame3.data[ 285] = 8'h10; frame3.valid[ 285] = 1'b1; frame3.error[ 285] = 1'b0;
        frame3.data[ 286] = 8'h11; frame3.valid[ 286] = 1'b1; frame3.error[ 286] = 1'b0;frame3.data[ 287] = 8'h12; frame3.valid[ 287] = 1'b1; frame3.error[ 287] = 1'b0;frame3.data[ 288] = 8'h13; frame3.valid[ 288] = 1'b1; frame3.error[ 288] = 1'b0;frame3.data[ 289] = 8'h14; frame3.valid[ 289] = 1'b1; frame3.error[ 289] = 1'b0;frame3.data[ 290] = 8'h15; frame3.valid[ 290] = 1'b1; frame3.error[ 290] = 1'b0;frame3.data[ 291] = 8'h16; frame3.valid[ 291] = 1'b1; frame3.error[ 291] = 1'b0;frame3.data[ 292] = 8'h17; frame3.valid[ 292] = 1'b1; frame3.error[ 292] = 1'b0;frame3.data[ 293] = 8'h18; frame3.valid[ 293] = 1'b1; frame3.error[ 293] = 1'b0;frame3.data[ 294] = 8'h19; frame3.valid[ 294] = 1'b1; frame3.error[ 294] = 1'b0;frame3.data[ 295] = 8'h1A; frame3.valid[ 295] = 1'b1; frame3.error[ 295] = 1'b0;frame3.data[ 296] = 8'h1B; frame3.valid[ 296] = 1'b1; frame3.error[ 296] = 1'b0;frame3.data[ 297] = 8'h1C; frame3.valid[ 297] = 1'b1; frame3.error[ 297] = 1'b0;frame3.data[ 298] = 8'h1D; frame3.valid[ 298] = 1'b1; frame3.error[ 298] = 1'b0;frame3.data[ 299] = 8'h1E; frame3.valid[ 299] = 1'b1; frame3.error[ 299] = 1'b0;frame3.data[ 300] = 8'h1F; frame3.valid[ 300] = 1'b1; frame3.error[ 300] = 1'b0;frame3.data[ 301] = 8'h20; frame3.valid[ 301] = 1'b1; frame3.error[ 301] = 1'b0;
        frame3.data[ 302] = 8'h21; frame3.valid[ 302] = 1'b1; frame3.error[ 302] = 1'b0;frame3.data[ 303] = 8'h22; frame3.valid[ 303] = 1'b1; frame3.error[ 303] = 1'b0;frame3.data[ 304] = 8'h23; frame3.valid[ 304] = 1'b1; frame3.error[ 304] = 1'b0;frame3.data[ 305] = 8'h24; frame3.valid[ 305] = 1'b1; frame3.error[ 305] = 1'b0;frame3.data[ 306] = 8'h25; frame3.valid[ 306] = 1'b1; frame3.error[ 306] = 1'b0;frame3.data[ 307] = 8'h26; frame3.valid[ 307] = 1'b1; frame3.error[ 307] = 1'b0;frame3.data[ 308] = 8'h27; frame3.valid[ 308] = 1'b1; frame3.error[ 308] = 1'b0;frame3.data[ 309] = 8'h28; frame3.valid[ 309] = 1'b1; frame3.error[ 309] = 1'b0;frame3.data[ 310] = 8'h29; frame3.valid[ 310] = 1'b1; frame3.error[ 310] = 1'b0;frame3.data[ 311] = 8'h2A; frame3.valid[ 311] = 1'b1; frame3.error[ 311] = 1'b0;frame3.data[ 312] = 8'h2B; frame3.valid[ 312] = 1'b1; frame3.error[ 312] = 1'b0;frame3.data[ 313] = 8'h2C; frame3.valid[ 313] = 1'b1; frame3.error[ 313] = 1'b0;frame3.data[ 314] = 8'h2D; frame3.valid[ 314] = 1'b1; frame3.error[ 314] = 1'b0;frame3.data[ 315] = 8'h2E; frame3.valid[ 315] = 1'b1; frame3.error[ 315] = 1'b0;frame3.data[ 316] = 8'h2F; frame3.valid[ 316] = 1'b1; frame3.error[ 316] = 1'b0;frame3.data[ 317] = 8'h30; frame3.valid[ 317] = 1'b1; frame3.error[ 317] = 1'b0;
        frame3.data[ 318] = 8'h31; frame3.valid[ 318] = 1'b1; frame3.error[ 318] = 1'b0;frame3.data[ 319] = 8'h32; frame3.valid[ 319] = 1'b1; frame3.error[ 319] = 1'b0;frame3.data[ 320] = 8'h33; frame3.valid[ 320] = 1'b1; frame3.error[ 320] = 1'b0;frame3.data[ 321] = 8'h34; frame3.valid[ 321] = 1'b1; frame3.error[ 321] = 1'b0;frame3.data[ 322] = 8'h35; frame3.valid[ 322] = 1'b1; frame3.error[ 322] = 1'b0;frame3.data[ 323] = 8'h36; frame3.valid[ 323] = 1'b1; frame3.error[ 323] = 1'b0;frame3.data[ 324] = 8'h37; frame3.valid[ 324] = 1'b1; frame3.error[ 324] = 1'b0;frame3.data[ 325] = 8'h38; frame3.valid[ 325] = 1'b1; frame3.error[ 325] = 1'b0;frame3.data[ 326] = 8'h39; frame3.valid[ 326] = 1'b1; frame3.error[ 326] = 1'b0;frame3.data[ 327] = 8'h3A; frame3.valid[ 327] = 1'b1; frame3.error[ 327] = 1'b0;frame3.data[ 328] = 8'h3B; frame3.valid[ 328] = 1'b1; frame3.error[ 328] = 1'b0;frame3.data[ 329] = 8'h3C; frame3.valid[ 329] = 1'b1; frame3.error[ 329] = 1'b0;frame3.data[ 330] = 8'h3D; frame3.valid[ 330] = 1'b1; frame3.error[ 330] = 1'b0;frame3.data[ 331] = 8'h3E; frame3.valid[ 331] = 1'b1; frame3.error[ 331] = 1'b0;frame3.data[ 332] = 8'h3F; frame3.valid[ 332] = 1'b1; frame3.error[ 332] = 1'b0;frame3.data[ 333] = 8'h40; frame3.valid[ 333] = 1'b1; frame3.error[ 333] = 1'b0;
        frame3.data[ 334] = 8'h41; frame3.valid[ 334] = 1'b1; frame3.error[ 334] = 1'b0;frame3.data[ 335] = 8'h42; frame3.valid[ 335] = 1'b1; frame3.error[ 335] = 1'b0;frame3.data[ 336] = 8'h43; frame3.valid[ 336] = 1'b1; frame3.error[ 336] = 1'b0;frame3.data[ 337] = 8'h44; frame3.valid[ 337] = 1'b1; frame3.error[ 337] = 1'b0;frame3.data[ 338] = 8'h45; frame3.valid[ 338] = 1'b1; frame3.error[ 338] = 1'b0;frame3.data[ 339] = 8'h46; frame3.valid[ 339] = 1'b1; frame3.error[ 339] = 1'b0;frame3.data[ 340] = 8'h47; frame3.valid[ 340] = 1'b1; frame3.error[ 340] = 1'b0;frame3.data[ 341] = 8'h48; frame3.valid[ 341] = 1'b1; frame3.error[ 341] = 1'b0;frame3.data[ 342] = 8'h49; frame3.valid[ 342] = 1'b1; frame3.error[ 342] = 1'b0;frame3.data[ 343] = 8'h4A; frame3.valid[ 343] = 1'b1; frame3.error[ 343] = 1'b0;frame3.data[ 344] = 8'h4B; frame3.valid[ 344] = 1'b1; frame3.error[ 344] = 1'b0;frame3.data[ 345] = 8'h4C; frame3.valid[ 345] = 1'b1; frame3.error[ 345] = 1'b0;frame3.data[ 346] = 8'h4D; frame3.valid[ 346] = 1'b1; frame3.error[ 346] = 1'b0;frame3.data[ 347] = 8'h4E; frame3.valid[ 347] = 1'b1; frame3.error[ 347] = 1'b0;frame3.data[ 348] = 8'h4F; frame3.valid[ 348] = 1'b1; frame3.error[ 348] = 1'b0;frame3.data[ 349] = 8'h50; frame3.valid[ 349] = 1'b1; frame3.error[ 349] = 1'b0;
        frame3.data[ 350] = 8'h51; frame3.valid[ 350] = 1'b1; frame3.error[ 350] = 1'b0;frame3.data[ 351] = 8'h52; frame3.valid[ 351] = 1'b1; frame3.error[ 351] = 1'b0;frame3.data[ 352] = 8'h53; frame3.valid[ 352] = 1'b1; frame3.error[ 352] = 1'b0;frame3.data[ 353] = 8'h54; frame3.valid[ 353] = 1'b1; frame3.error[ 353] = 1'b0;frame3.data[ 354] = 8'h55; frame3.valid[ 354] = 1'b1; frame3.error[ 354] = 1'b0;frame3.data[ 355] = 8'h56; frame3.valid[ 355] = 1'b1; frame3.error[ 355] = 1'b0;frame3.data[ 356] = 8'h57; frame3.valid[ 356] = 1'b1; frame3.error[ 356] = 1'b0;frame3.data[ 357] = 8'h58; frame3.valid[ 357] = 1'b1; frame3.error[ 357] = 1'b0;frame3.data[ 358] = 8'h59; frame3.valid[ 358] = 1'b1; frame3.error[ 358] = 1'b0;frame3.data[ 359] = 8'h5A; frame3.valid[ 359] = 1'b1; frame3.error[ 359] = 1'b0;frame3.data[ 360] = 8'h5B; frame3.valid[ 360] = 1'b1; frame3.error[ 360] = 1'b0;frame3.data[ 361] = 8'h5C; frame3.valid[ 361] = 1'b1; frame3.error[ 361] = 1'b0;frame3.data[ 362] = 8'h5D; frame3.valid[ 362] = 1'b1; frame3.error[ 362] = 1'b0;frame3.data[ 363] = 8'h5E; frame3.valid[ 363] = 1'b1; frame3.error[ 363] = 1'b0;frame3.data[ 364] = 8'h5F; frame3.valid[ 364] = 1'b1; frame3.error[ 364] = 1'b0;frame3.data[ 365] = 8'h60; frame3.valid[ 365] = 1'b1; frame3.error[ 365] = 1'b0;
        frame3.data[ 366] = 8'h61; frame3.valid[ 366] = 1'b1; frame3.error[ 366] = 1'b0;frame3.data[ 367] = 8'h62; frame3.valid[ 367] = 1'b1; frame3.error[ 367] = 1'b0;frame3.data[ 368] = 8'h63; frame3.valid[ 368] = 1'b1; frame3.error[ 368] = 1'b0;frame3.data[ 369] = 8'h64; frame3.valid[ 369] = 1'b1; frame3.error[ 369] = 1'b0;frame3.data[ 370] = 8'h65; frame3.valid[ 370] = 1'b1; frame3.error[ 370] = 1'b0;frame3.data[ 371] = 8'h66; frame3.valid[ 371] = 1'b1; frame3.error[ 371] = 1'b0;frame3.data[ 372] = 8'h67; frame3.valid[ 372] = 1'b1; frame3.error[ 372] = 1'b0;frame3.data[ 373] = 8'h68; frame3.valid[ 373] = 1'b1; frame3.error[ 373] = 1'b0;frame3.data[ 374] = 8'h69; frame3.valid[ 374] = 1'b1; frame3.error[ 374] = 1'b0;frame3.data[ 375] = 8'h6A; frame3.valid[ 375] = 1'b1; frame3.error[ 375] = 1'b0;frame3.data[ 376] = 8'h6B; frame3.valid[ 376] = 1'b1; frame3.error[ 376] = 1'b0;frame3.data[ 377] = 8'h6C; frame3.valid[ 377] = 1'b1; frame3.error[ 377] = 1'b0;frame3.data[ 378] = 8'h6D; frame3.valid[ 378] = 1'b1; frame3.error[ 378] = 1'b0;frame3.data[ 379] = 8'h6E; frame3.valid[ 379] = 1'b1; frame3.error[ 379] = 1'b0;frame3.data[ 380] = 8'h6F; frame3.valid[ 380] = 1'b1; frame3.error[ 380] = 1'b0;frame3.data[ 381] = 8'h70; frame3.valid[ 381] = 1'b1; frame3.error[ 381] = 1'b0;
        frame3.data[ 382] = 8'h71; frame3.valid[ 382] = 1'b1; frame3.error[ 382] = 1'b0;frame3.data[ 383] = 8'h72; frame3.valid[ 383] = 1'b1; frame3.error[ 383] = 1'b0;frame3.data[ 384] = 8'h73; frame3.valid[ 384] = 1'b1; frame3.error[ 384] = 1'b0;frame3.data[ 385] = 8'h74; frame3.valid[ 385] = 1'b1; frame3.error[ 385] = 1'b0;frame3.data[ 386] = 8'h75; frame3.valid[ 386] = 1'b1; frame3.error[ 386] = 1'b0;frame3.data[ 387] = 8'h76; frame3.valid[ 387] = 1'b1; frame3.error[ 387] = 1'b0;frame3.data[ 388] = 8'h77; frame3.valid[ 388] = 1'b1; frame3.error[ 388] = 1'b0;frame3.data[ 389] = 8'h78; frame3.valid[ 389] = 1'b1; frame3.error[ 389] = 1'b0;frame3.data[ 390] = 8'h79; frame3.valid[ 390] = 1'b1; frame3.error[ 390] = 1'b0;frame3.data[ 391] = 8'h7A; frame3.valid[ 391] = 1'b1; frame3.error[ 391] = 1'b0;frame3.data[ 392] = 8'h7B; frame3.valid[ 392] = 1'b1; frame3.error[ 392] = 1'b0;frame3.data[ 393] = 8'h7C; frame3.valid[ 393] = 1'b1; frame3.error[ 393] = 1'b0;frame3.data[ 394] = 8'h7D; frame3.valid[ 394] = 1'b1; frame3.error[ 394] = 1'b0;frame3.data[ 395] = 8'h7E; frame3.valid[ 395] = 1'b1; frame3.error[ 395] = 1'b0;frame3.data[ 396] = 8'h7F; frame3.valid[ 396] = 1'b1; frame3.error[ 396] = 1'b0;frame3.data[ 397] = 8'h80; frame3.valid[ 397] = 1'b1; frame3.error[ 397] = 1'b0;
        frame3.data[ 398] = 8'h81; frame3.valid[ 398] = 1'b1; frame3.error[ 398] = 1'b0;frame3.data[ 399] = 8'h82; frame3.valid[ 399] = 1'b1; frame3.error[ 399] = 1'b0;frame3.data[ 400] = 8'h83; frame3.valid[ 400] = 1'b1; frame3.error[ 400] = 1'b0;frame3.data[ 401] = 8'h84; frame3.valid[ 401] = 1'b1; frame3.error[ 401] = 1'b0;frame3.data[ 402] = 8'h85; frame3.valid[ 402] = 1'b1; frame3.error[ 402] = 1'b0;frame3.data[ 403] = 8'h86; frame3.valid[ 403] = 1'b1; frame3.error[ 403] = 1'b0;frame3.data[ 404] = 8'h87; frame3.valid[ 404] = 1'b1; frame3.error[ 404] = 1'b0;frame3.data[ 405] = 8'h88; frame3.valid[ 405] = 1'b1; frame3.error[ 405] = 1'b0;frame3.data[ 406] = 8'h89; frame3.valid[ 406] = 1'b1; frame3.error[ 406] = 1'b0;frame3.data[ 407] = 8'h8A; frame3.valid[ 407] = 1'b1; frame3.error[ 407] = 1'b0;frame3.data[ 408] = 8'h8B; frame3.valid[ 408] = 1'b1; frame3.error[ 408] = 1'b0;frame3.data[ 409] = 8'h8C; frame3.valid[ 409] = 1'b1; frame3.error[ 409] = 1'b0;frame3.data[ 410] = 8'h8D; frame3.valid[ 410] = 1'b1; frame3.error[ 410] = 1'b0;frame3.data[ 411] = 8'h8E; frame3.valid[ 411] = 1'b1; frame3.error[ 411] = 1'b0;frame3.data[ 412] = 8'h8F; frame3.valid[ 412] = 1'b1; frame3.error[ 412] = 1'b0;frame3.data[ 413] = 8'h90; frame3.valid[ 413] = 1'b1; frame3.error[ 413] = 1'b0;
        frame3.data[ 414] = 8'h91; frame3.valid[ 414] = 1'b1; frame3.error[ 414] = 1'b0;frame3.data[ 415] = 8'h92; frame3.valid[ 415] = 1'b1; frame3.error[ 415] = 1'b0;frame3.data[ 416] = 8'h93; frame3.valid[ 416] = 1'b1; frame3.error[ 416] = 1'b0;frame3.data[ 417] = 8'h94; frame3.valid[ 417] = 1'b1; frame3.error[ 417] = 1'b0;frame3.data[ 418] = 8'h95; frame3.valid[ 418] = 1'b1; frame3.error[ 418] = 1'b0;frame3.data[ 419] = 8'h96; frame3.valid[ 419] = 1'b1; frame3.error[ 419] = 1'b0;frame3.data[ 420] = 8'h97; frame3.valid[ 420] = 1'b1; frame3.error[ 420] = 1'b0;frame3.data[ 421] = 8'h98; frame3.valid[ 421] = 1'b1; frame3.error[ 421] = 1'b0;frame3.data[ 422] = 8'h99; frame3.valid[ 422] = 1'b1; frame3.error[ 422] = 1'b0;frame3.data[ 423] = 8'h9A; frame3.valid[ 423] = 1'b1; frame3.error[ 423] = 1'b0;frame3.data[ 424] = 8'h9B; frame3.valid[ 424] = 1'b1; frame3.error[ 424] = 1'b0;frame3.data[ 425] = 8'h9C; frame3.valid[ 425] = 1'b1; frame3.error[ 425] = 1'b0;frame3.data[ 426] = 8'h9D; frame3.valid[ 426] = 1'b1; frame3.error[ 426] = 1'b0;frame3.data[ 427] = 8'h9E; frame3.valid[ 427] = 1'b1; frame3.error[ 427] = 1'b0;frame3.data[ 428] = 8'h9F; frame3.valid[ 428] = 1'b1; frame3.error[ 428] = 1'b0;frame3.data[ 429] = 8'hA0; frame3.valid[ 429] = 1'b1; frame3.error[ 429] = 1'b0;
        frame3.data[ 430] = 8'hA1; frame3.valid[ 430] = 1'b1; frame3.error[ 430] = 1'b0;frame3.data[ 431] = 8'hA2; frame3.valid[ 431] = 1'b1; frame3.error[ 431] = 1'b0;frame3.data[ 432] = 8'hA3; frame3.valid[ 432] = 1'b1; frame3.error[ 432] = 1'b0;frame3.data[ 433] = 8'hA4; frame3.valid[ 433] = 1'b1; frame3.error[ 433] = 1'b0;frame3.data[ 434] = 8'hA5; frame3.valid[ 434] = 1'b1; frame3.error[ 434] = 1'b0;frame3.data[ 435] = 8'hA6; frame3.valid[ 435] = 1'b1; frame3.error[ 435] = 1'b0;frame3.data[ 436] = 8'hA7; frame3.valid[ 436] = 1'b1; frame3.error[ 436] = 1'b0;frame3.data[ 437] = 8'hA8; frame3.valid[ 437] = 1'b1; frame3.error[ 437] = 1'b0;frame3.data[ 438] = 8'hA9; frame3.valid[ 438] = 1'b1; frame3.error[ 438] = 1'b0;frame3.data[ 439] = 8'hAA; frame3.valid[ 439] = 1'b1; frame3.error[ 439] = 1'b0;frame3.data[ 440] = 8'hAB; frame3.valid[ 440] = 1'b1; frame3.error[ 440] = 1'b0;frame3.data[ 441] = 8'hAC; frame3.valid[ 441] = 1'b1; frame3.error[ 441] = 1'b0;frame3.data[ 442] = 8'hAD; frame3.valid[ 442] = 1'b1; frame3.error[ 442] = 1'b0;frame3.data[ 443] = 8'hAE; frame3.valid[ 443] = 1'b1; frame3.error[ 443] = 1'b0;frame3.data[ 444] = 8'hAF; frame3.valid[ 444] = 1'b1; frame3.error[ 444] = 1'b0;frame3.data[ 445] = 8'hB0; frame3.valid[ 445] = 1'b1; frame3.error[ 445] = 1'b0;
        frame3.data[ 446] = 8'hB1; frame3.valid[ 446] = 1'b1; frame3.error[ 446] = 1'b0;frame3.data[ 447] = 8'hB2; frame3.valid[ 447] = 1'b1; frame3.error[ 447] = 1'b0;frame3.data[ 448] = 8'hB3; frame3.valid[ 448] = 1'b1; frame3.error[ 448] = 1'b0;frame3.data[ 449] = 8'hB4; frame3.valid[ 449] = 1'b1; frame3.error[ 449] = 1'b0;frame3.data[ 450] = 8'hB5; frame3.valid[ 450] = 1'b1; frame3.error[ 450] = 1'b0;frame3.data[ 451] = 8'hB6; frame3.valid[ 451] = 1'b1; frame3.error[ 451] = 1'b0;frame3.data[ 452] = 8'hB7; frame3.valid[ 452] = 1'b1; frame3.error[ 452] = 1'b0;frame3.data[ 453] = 8'hB8; frame3.valid[ 453] = 1'b1; frame3.error[ 453] = 1'b0;frame3.data[ 454] = 8'hB9; frame3.valid[ 454] = 1'b1; frame3.error[ 454] = 1'b0;frame3.data[ 455] = 8'hBA; frame3.valid[ 455] = 1'b1; frame3.error[ 455] = 1'b0;frame3.data[ 456] = 8'hBB; frame3.valid[ 456] = 1'b1; frame3.error[ 456] = 1'b0;frame3.data[ 457] = 8'hBC; frame3.valid[ 457] = 1'b1; frame3.error[ 457] = 1'b0;frame3.data[ 458] = 8'hBD; frame3.valid[ 458] = 1'b1; frame3.error[ 458] = 1'b0;frame3.data[ 459] = 8'hBE; frame3.valid[ 459] = 1'b1; frame3.error[ 459] = 1'b0;frame3.data[ 460] = 8'hBF; frame3.valid[ 460] = 1'b1; frame3.error[ 460] = 1'b0;frame3.data[ 461] = 8'hC0; frame3.valid[ 461] = 1'b1; frame3.error[ 461] = 1'b0;
        frame3.data[ 462] = 8'hC1; frame3.valid[ 462] = 1'b1; frame3.error[ 462] = 1'b0;frame3.data[ 463] = 8'hC2; frame3.valid[ 463] = 1'b1; frame3.error[ 463] = 1'b0;frame3.data[ 464] = 8'hC3; frame3.valid[ 464] = 1'b1; frame3.error[ 464] = 1'b0;frame3.data[ 465] = 8'hC4; frame3.valid[ 465] = 1'b1; frame3.error[ 465] = 1'b0;frame3.data[ 466] = 8'hC5; frame3.valid[ 466] = 1'b1; frame3.error[ 466] = 1'b0;frame3.data[ 467] = 8'hC6; frame3.valid[ 467] = 1'b1; frame3.error[ 467] = 1'b0;frame3.data[ 468] = 8'hC7; frame3.valid[ 468] = 1'b1; frame3.error[ 468] = 1'b0;frame3.data[ 469] = 8'hC8; frame3.valid[ 469] = 1'b1; frame3.error[ 469] = 1'b0;frame3.data[ 470] = 8'hC9; frame3.valid[ 470] = 1'b1; frame3.error[ 470] = 1'b0;frame3.data[ 471] = 8'hCA; frame3.valid[ 471] = 1'b1; frame3.error[ 471] = 1'b0;frame3.data[ 472] = 8'hCB; frame3.valid[ 472] = 1'b1; frame3.error[ 472] = 1'b0;frame3.data[ 473] = 8'hCC; frame3.valid[ 473] = 1'b1; frame3.error[ 473] = 1'b0;frame3.data[ 474] = 8'hCD; frame3.valid[ 474] = 1'b1; frame3.error[ 474] = 1'b0;frame3.data[ 475] = 8'hCE; frame3.valid[ 475] = 1'b1; frame3.error[ 475] = 1'b0;frame3.data[ 476] = 8'hCF; frame3.valid[ 476] = 1'b1; frame3.error[ 476] = 1'b0;frame3.data[ 477] = 8'hD0; frame3.valid[ 477] = 1'b1; frame3.error[ 477] = 1'b0;
        frame3.data[ 478] = 8'hD1; frame3.valid[ 478] = 1'b1; frame3.error[ 478] = 1'b0;frame3.data[ 479] = 8'hD2; frame3.valid[ 479] = 1'b1; frame3.error[ 479] = 1'b0;frame3.data[ 480] = 8'hD3; frame3.valid[ 480] = 1'b1; frame3.error[ 480] = 1'b0;frame3.data[ 481] = 8'hD4; frame3.valid[ 481] = 1'b1; frame3.error[ 481] = 1'b0;frame3.data[ 482] = 8'hD5; frame3.valid[ 482] = 1'b1; frame3.error[ 482] = 1'b0;frame3.data[ 483] = 8'hD6; frame3.valid[ 483] = 1'b1; frame3.error[ 483] = 1'b0;frame3.data[ 484] = 8'hD7; frame3.valid[ 484] = 1'b1; frame3.error[ 484] = 1'b0;frame3.data[ 485] = 8'hD8; frame3.valid[ 485] = 1'b1; frame3.error[ 485] = 1'b0;frame3.data[ 486] = 8'hD9; frame3.valid[ 486] = 1'b1; frame3.error[ 486] = 1'b0;frame3.data[ 487] = 8'hDA; frame3.valid[ 487] = 1'b1; frame3.error[ 487] = 1'b0;frame3.data[ 488] = 8'hDB; frame3.valid[ 488] = 1'b1; frame3.error[ 488] = 1'b0;frame3.data[ 489] = 8'hDC; frame3.valid[ 489] = 1'b1; frame3.error[ 489] = 1'b0;frame3.data[ 490] = 8'hDD; frame3.valid[ 490] = 1'b1; frame3.error[ 490] = 1'b0;frame3.data[ 491] = 8'hDE; frame3.valid[ 491] = 1'b1; frame3.error[ 491] = 1'b0;frame3.data[ 492] = 8'hDF; frame3.valid[ 492] = 1'b1; frame3.error[ 492] = 1'b0;frame3.data[ 493] = 8'hE0; frame3.valid[ 493] = 1'b1; frame3.error[ 493] = 1'b0;
        frame3.data[ 494] = 8'hE1; frame3.valid[ 494] = 1'b1; frame3.error[ 494] = 1'b0;frame3.data[ 495] = 8'hE2; frame3.valid[ 495] = 1'b1; frame3.error[ 495] = 1'b0;frame3.data[ 496] = 8'hE3; frame3.valid[ 496] = 1'b1; frame3.error[ 496] = 1'b0;frame3.data[ 497] = 8'hE4; frame3.valid[ 497] = 1'b1; frame3.error[ 497] = 1'b0;frame3.data[ 498] = 8'hE5; frame3.valid[ 498] = 1'b1; frame3.error[ 498] = 1'b0;frame3.data[ 499] = 8'hE6; frame3.valid[ 499] = 1'b1; frame3.error[ 499] = 1'b0;frame3.data[ 500] = 8'hE7; frame3.valid[ 500] = 1'b1; frame3.error[ 500] = 1'b0;frame3.data[ 501] = 8'hE8; frame3.valid[ 501] = 1'b1; frame3.error[ 501] = 1'b0;frame3.data[ 502] = 8'hE9; frame3.valid[ 502] = 1'b1; frame3.error[ 502] = 1'b0;frame3.data[ 503] = 8'hEA; frame3.valid[ 503] = 1'b1; frame3.error[ 503] = 1'b0;frame3.data[ 504] = 8'hEB; frame3.valid[ 504] = 1'b1; frame3.error[ 504] = 1'b0;frame3.data[ 505] = 8'hEC; frame3.valid[ 505] = 1'b1; frame3.error[ 505] = 1'b0;frame3.data[ 506] = 8'hED; frame3.valid[ 506] = 1'b1; frame3.error[ 506] = 1'b0;frame3.data[ 507] = 8'hEE; frame3.valid[ 507] = 1'b1; frame3.error[ 507] = 1'b0;frame3.data[ 508] = 8'hEF; frame3.valid[ 508] = 1'b1; frame3.error[ 508] = 1'b0;frame3.data[ 509] = 8'hF0; frame3.valid[ 509] = 1'b1; frame3.error[ 509] = 1'b0;
        frame3.data[ 510] = 8'hF1; frame3.valid[ 510] = 1'b1; frame3.error[ 510] = 1'b0;frame3.data[ 511] = 8'hF2; frame3.valid[ 511] = 1'b1; frame3.error[ 511] = 1'b0;frame3.data[ 512] = 8'hF3; frame3.valid[ 512] = 1'b1; frame3.error[ 512] = 1'b0;frame3.data[ 513] = 8'hF4; frame3.valid[ 513] = 1'b1; frame3.error[ 513] = 1'b0;frame3.data[ 514] = 8'hF5; frame3.valid[ 514] = 1'b1; frame3.error[ 514] = 1'b0;frame3.data[ 515] = 8'hF6; frame3.valid[ 515] = 1'b1; frame3.error[ 515] = 1'b0;frame3.data[ 516] = 8'hF7; frame3.valid[ 516] = 1'b1; frame3.error[ 516] = 1'b0;frame3.data[ 517] = 8'hF8; frame3.valid[ 517] = 1'b1; frame3.error[ 517] = 1'b0;frame3.data[ 518] = 8'hF9; frame3.valid[ 518] = 1'b1; frame3.error[ 518] = 1'b0;frame3.data[ 519] = 8'hFA; frame3.valid[ 519] = 1'b1; frame3.error[ 519] = 1'b0;frame3.data[ 520] = 8'hFB; frame3.valid[ 520] = 1'b1; frame3.error[ 520] = 1'b0;frame3.data[ 521] = 8'hFC; frame3.valid[ 521] = 1'b1; frame3.error[ 521] = 1'b0;frame3.data[ 522] = 8'hFD; frame3.valid[ 522] = 1'b1; frame3.error[ 522] = 1'b0;frame3.data[ 523] = 8'hFE; frame3.valid[ 523] = 1'b1; frame3.error[ 523] = 1'b0;frame3.data[ 524] = 8'h00; frame3.valid[ 524] = 1'b1; frame3.error[ 524] = 1'b0;frame3.data[ 525] = 8'h01; frame3.valid[ 525] = 1'b1; frame3.error[ 525] = 1'b0;
        frame3.data[ 526] = 8'h02; frame3.valid[ 526] = 1'b1; frame3.error[ 526] = 1'b0;frame3.data[ 527] = 8'h03; frame3.valid[ 527] = 1'b1; frame3.error[ 527] = 1'b0;frame3.data[ 528] = 8'h04; frame3.valid[ 528] = 1'b1; frame3.error[ 528] = 1'b0;frame3.data[ 529] = 8'h05; frame3.valid[ 529] = 1'b1; frame3.error[ 529] = 1'b0;frame3.data[ 530] = 8'h06; frame3.valid[ 530] = 1'b1; frame3.error[ 530] = 1'b0;frame3.data[ 531] = 8'h07; frame3.valid[ 531] = 1'b1; frame3.error[ 531] = 1'b0;frame3.data[ 532] = 8'h08; frame3.valid[ 532] = 1'b1; frame3.error[ 532] = 1'b0;frame3.data[ 533] = 8'h09; frame3.valid[ 533] = 1'b1; frame3.error[ 533] = 1'b0;frame3.data[ 534] = 8'h0A; frame3.valid[ 534] = 1'b1; frame3.error[ 534] = 1'b0;frame3.data[ 535] = 8'h0B; frame3.valid[ 535] = 1'b1; frame3.error[ 535] = 1'b0;frame3.data[ 536] = 8'h0C; frame3.valid[ 536] = 1'b1; frame3.error[ 536] = 1'b0;frame3.data[ 537] = 8'h0D; frame3.valid[ 537] = 1'b1; frame3.error[ 537] = 1'b0;frame3.data[ 538] = 8'h0E; frame3.valid[ 538] = 1'b1; frame3.error[ 538] = 1'b0;frame3.data[ 539] = 8'h0F; frame3.valid[ 539] = 1'b1; frame3.error[ 539] = 1'b0;frame3.data[ 540] = 8'h10; frame3.valid[ 540] = 1'b1; frame3.error[ 540] = 1'b0;frame3.data[ 541] = 8'h11; frame3.valid[ 541] = 1'b1; frame3.error[ 541] = 1'b0;
        frame3.data[ 542] = 8'h12; frame3.valid[ 542] = 1'b1; frame3.error[ 542] = 1'b0;frame3.data[ 543] = 8'h13; frame3.valid[ 543] = 1'b1; frame3.error[ 543] = 1'b0;frame3.data[ 544] = 8'h14; frame3.valid[ 544] = 1'b1; frame3.error[ 544] = 1'b0;frame3.data[ 545] = 8'h15; frame3.valid[ 545] = 1'b1; frame3.error[ 545] = 1'b0;frame3.data[ 546] = 8'h16; frame3.valid[ 546] = 1'b1; frame3.error[ 546] = 1'b0;frame3.data[ 547] = 8'h17; frame3.valid[ 547] = 1'b1; frame3.error[ 547] = 1'b0;frame3.data[ 548] = 8'h18; frame3.valid[ 548] = 1'b1; frame3.error[ 548] = 1'b0;frame3.data[ 549] = 8'h19; frame3.valid[ 549] = 1'b1; frame3.error[ 549] = 1'b0;frame3.data[ 550] = 8'h1A; frame3.valid[ 550] = 1'b1; frame3.error[ 550] = 1'b0;frame3.data[ 551] = 8'h1B; frame3.valid[ 551] = 1'b1; frame3.error[ 551] = 1'b0;frame3.data[ 552] = 8'h1C; frame3.valid[ 552] = 1'b1; frame3.error[ 552] = 1'b0;frame3.data[ 553] = 8'h1D; frame3.valid[ 553] = 1'b1; frame3.error[ 553] = 1'b0;frame3.data[ 554] = 8'h1E; frame3.valid[ 554] = 1'b1; frame3.error[ 554] = 1'b0;frame3.data[ 555] = 8'h1F; frame3.valid[ 555] = 1'b1; frame3.error[ 555] = 1'b0;frame3.data[ 556] = 8'h20; frame3.valid[ 556] = 1'b1; frame3.error[ 556] = 1'b0;frame3.data[ 557] = 8'h21; frame3.valid[ 557] = 1'b1; frame3.error[ 557] = 1'b0;
        frame3.data[ 558] = 8'h22; frame3.valid[ 558] = 1'b1; frame3.error[ 558] = 1'b0;frame3.data[ 559] = 8'h23; frame3.valid[ 559] = 1'b1; frame3.error[ 559] = 1'b0;frame3.data[ 560] = 8'h24; frame3.valid[ 560] = 1'b1; frame3.error[ 560] = 1'b0;frame3.data[ 561] = 8'h25; frame3.valid[ 561] = 1'b1; frame3.error[ 561] = 1'b0;frame3.data[ 562] = 8'h26; frame3.valid[ 562] = 1'b1; frame3.error[ 562] = 1'b0;frame3.data[ 563] = 8'h27; frame3.valid[ 563] = 1'b1; frame3.error[ 563] = 1'b0;frame3.data[ 564] = 8'h28; frame3.valid[ 564] = 1'b1; frame3.error[ 564] = 1'b0;frame3.data[ 565] = 8'h29; frame3.valid[ 565] = 1'b1; frame3.error[ 565] = 1'b0;frame3.data[ 566] = 8'h2A; frame3.valid[ 566] = 1'b1; frame3.error[ 566] = 1'b0;frame3.data[ 567] = 8'h2B; frame3.valid[ 567] = 1'b1; frame3.error[ 567] = 1'b0;frame3.data[ 568] = 8'h2C; frame3.valid[ 568] = 1'b1; frame3.error[ 568] = 1'b0;frame3.data[ 569] = 8'h2D; frame3.valid[ 569] = 1'b1; frame3.error[ 569] = 1'b0;frame3.data[ 570] = 8'h2E; frame3.valid[ 570] = 1'b1; frame3.error[ 570] = 1'b0;frame3.data[ 571] = 8'h2F; frame3.valid[ 571] = 1'b1; frame3.error[ 571] = 1'b0;frame3.data[ 572] = 8'h30; frame3.valid[ 572] = 1'b1; frame3.error[ 572] = 1'b0;frame3.data[ 573] = 8'h31; frame3.valid[ 573] = 1'b1; frame3.error[ 573] = 1'b0;
        frame3.data[ 574] = 8'h32; frame3.valid[ 574] = 1'b1; frame3.error[ 574] = 1'b0;frame3.data[ 575] = 8'h33; frame3.valid[ 575] = 1'b1; frame3.error[ 575] = 1'b0;frame3.data[ 576] = 8'h34; frame3.valid[ 576] = 1'b1; frame3.error[ 576] = 1'b0;frame3.data[ 577] = 8'h35; frame3.valid[ 577] = 1'b1; frame3.error[ 577] = 1'b0;frame3.data[ 578] = 8'h36; frame3.valid[ 578] = 1'b1; frame3.error[ 578] = 1'b0;frame3.data[ 579] = 8'h37; frame3.valid[ 579] = 1'b1; frame3.error[ 579] = 1'b0;frame3.data[ 580] = 8'h38; frame3.valid[ 580] = 1'b1; frame3.error[ 580] = 1'b0;frame3.data[ 581] = 8'h39; frame3.valid[ 581] = 1'b1; frame3.error[ 581] = 1'b0;frame3.data[ 582] = 8'h3A; frame3.valid[ 582] = 1'b1; frame3.error[ 582] = 1'b0;frame3.data[ 583] = 8'h3B; frame3.valid[ 583] = 1'b1; frame3.error[ 583] = 1'b0;frame3.data[ 584] = 8'h3C; frame3.valid[ 584] = 1'b1; frame3.error[ 584] = 1'b0;frame3.data[ 585] = 8'h3D; frame3.valid[ 585] = 1'b1; frame3.error[ 585] = 1'b0;frame3.data[ 586] = 8'h3E; frame3.valid[ 586] = 1'b1; frame3.error[ 586] = 1'b0;frame3.data[ 587] = 8'h3F; frame3.valid[ 587] = 1'b1; frame3.error[ 587] = 1'b0;frame3.data[ 588] = 8'h40; frame3.valid[ 588] = 1'b1; frame3.error[ 588] = 1'b0;frame3.data[ 589] = 8'h41; frame3.valid[ 589] = 1'b1; frame3.error[ 589] = 1'b0;
        frame3.data[ 590] = 8'h42; frame3.valid[ 590] = 1'b1; frame3.error[ 590] = 1'b0;frame3.data[ 591] = 8'h43; frame3.valid[ 591] = 1'b1; frame3.error[ 591] = 1'b0;frame3.data[ 592] = 8'h44; frame3.valid[ 592] = 1'b1; frame3.error[ 592] = 1'b0;frame3.data[ 593] = 8'h45; frame3.valid[ 593] = 1'b1; frame3.error[ 593] = 1'b0;frame3.data[ 594] = 8'h46; frame3.valid[ 594] = 1'b1; frame3.error[ 594] = 1'b0;frame3.data[ 595] = 8'h47; frame3.valid[ 595] = 1'b1; frame3.error[ 595] = 1'b0;frame3.data[ 596] = 8'h48; frame3.valid[ 596] = 1'b1; frame3.error[ 596] = 1'b0;frame3.data[ 597] = 8'h49; frame3.valid[ 597] = 1'b1; frame3.error[ 597] = 1'b0;frame3.data[ 598] = 8'h4A; frame3.valid[ 598] = 1'b1; frame3.error[ 598] = 1'b0;frame3.data[ 599] = 8'h4B; frame3.valid[ 599] = 1'b1; frame3.error[ 599] = 1'b0;frame3.data[ 600] = 8'h4C; frame3.valid[ 600] = 1'b1; frame3.error[ 600] = 1'b0;frame3.data[ 601] = 8'h4D; frame3.valid[ 601] = 1'b1; frame3.error[ 601] = 1'b0;frame3.data[ 602] = 8'h4E; frame3.valid[ 602] = 1'b1; frame3.error[ 602] = 1'b0;frame3.data[ 603] = 8'h4F; frame3.valid[ 603] = 1'b1; frame3.error[ 603] = 1'b0;frame3.data[ 604] = 8'h50; frame3.valid[ 604] = 1'b1; frame3.error[ 604] = 1'b0;frame3.data[ 605] = 8'h51; frame3.valid[ 605] = 1'b1; frame3.error[ 605] = 1'b0;
        frame3.data[ 606] = 8'h52; frame3.valid[ 606] = 1'b1; frame3.error[ 606] = 1'b0;frame3.data[ 607] = 8'h53; frame3.valid[ 607] = 1'b1; frame3.error[ 607] = 1'b0;frame3.data[ 608] = 8'h54; frame3.valid[ 608] = 1'b1; frame3.error[ 608] = 1'b0;frame3.data[ 609] = 8'h55; frame3.valid[ 609] = 1'b1; frame3.error[ 609] = 1'b0;frame3.data[ 610] = 8'h56; frame3.valid[ 610] = 1'b1; frame3.error[ 610] = 1'b0;frame3.data[ 611] = 8'h57; frame3.valid[ 611] = 1'b1; frame3.error[ 611] = 1'b0;frame3.data[ 612] = 8'h58; frame3.valid[ 612] = 1'b1; frame3.error[ 612] = 1'b0;frame3.data[ 613] = 8'h59; frame3.valid[ 613] = 1'b1; frame3.error[ 613] = 1'b0;frame3.data[ 614] = 8'h5A; frame3.valid[ 614] = 1'b1; frame3.error[ 614] = 1'b0;frame3.data[ 615] = 8'h5B; frame3.valid[ 615] = 1'b1; frame3.error[ 615] = 1'b0;frame3.data[ 616] = 8'h5C; frame3.valid[ 616] = 1'b1; frame3.error[ 616] = 1'b0;frame3.data[ 617] = 8'h5D; frame3.valid[ 617] = 1'b1; frame3.error[ 617] = 1'b0;frame3.data[ 618] = 8'h5E; frame3.valid[ 618] = 1'b1; frame3.error[ 618] = 1'b0;frame3.data[ 619] = 8'h5F; frame3.valid[ 619] = 1'b1; frame3.error[ 619] = 1'b0;frame3.data[ 620] = 8'h60; frame3.valid[ 620] = 1'b1; frame3.error[ 620] = 1'b0;frame3.data[ 621] = 8'h61; frame3.valid[ 621] = 1'b1; frame3.error[ 621] = 1'b0;
        frame3.data[ 622] = 8'h62; frame3.valid[ 622] = 1'b1; frame3.error[ 622] = 1'b0;frame3.data[ 623] = 8'h63; frame3.valid[ 623] = 1'b1; frame3.error[ 623] = 1'b0;frame3.data[ 624] = 8'h64; frame3.valid[ 624] = 1'b1; frame3.error[ 624] = 1'b0;frame3.data[ 625] = 8'h65; frame3.valid[ 625] = 1'b1; frame3.error[ 625] = 1'b0;frame3.data[ 626] = 8'h66; frame3.valid[ 626] = 1'b1; frame3.error[ 626] = 1'b0;frame3.data[ 627] = 8'h67; frame3.valid[ 627] = 1'b1; frame3.error[ 627] = 1'b0;frame3.data[ 628] = 8'h68; frame3.valid[ 628] = 1'b1; frame3.error[ 628] = 1'b0;frame3.data[ 629] = 8'h69; frame3.valid[ 629] = 1'b1; frame3.error[ 629] = 1'b0;frame3.data[ 630] = 8'h6A; frame3.valid[ 630] = 1'b1; frame3.error[ 630] = 1'b0;frame3.data[ 631] = 8'h6B; frame3.valid[ 631] = 1'b1; frame3.error[ 631] = 1'b0;frame3.data[ 632] = 8'h6C; frame3.valid[ 632] = 1'b1; frame3.error[ 632] = 1'b0;frame3.data[ 633] = 8'h6D; frame3.valid[ 633] = 1'b1; frame3.error[ 633] = 1'b0;frame3.data[ 634] = 8'h6E; frame3.valid[ 634] = 1'b1; frame3.error[ 634] = 1'b0;frame3.data[ 635] = 8'h6F; frame3.valid[ 635] = 1'b1; frame3.error[ 635] = 1'b0;frame3.data[ 636] = 8'h70; frame3.valid[ 636] = 1'b1; frame3.error[ 636] = 1'b0;frame3.data[ 637] = 8'h71; frame3.valid[ 637] = 1'b1; frame3.error[ 637] = 1'b0;
        frame3.data[ 638] = 8'h72; frame3.valid[ 638] = 1'b1; frame3.error[ 638] = 1'b0;frame3.data[ 639] = 8'h73; frame3.valid[ 639] = 1'b1; frame3.error[ 639] = 1'b0;frame3.data[ 640] = 8'h74; frame3.valid[ 640] = 1'b1; frame3.error[ 640] = 1'b0;frame3.data[ 641] = 8'h75; frame3.valid[ 641] = 1'b1; frame3.error[ 641] = 1'b0;frame3.data[ 642] = 8'h76; frame3.valid[ 642] = 1'b1; frame3.error[ 642] = 1'b0;frame3.data[ 643] = 8'h77; frame3.valid[ 643] = 1'b1; frame3.error[ 643] = 1'b0;frame3.data[ 644] = 8'h78; frame3.valid[ 644] = 1'b1; frame3.error[ 644] = 1'b0;frame3.data[ 645] = 8'h79; frame3.valid[ 645] = 1'b1; frame3.error[ 645] = 1'b0;frame3.data[ 646] = 8'h7A; frame3.valid[ 646] = 1'b1; frame3.error[ 646] = 1'b0;frame3.data[ 647] = 8'h7B; frame3.valid[ 647] = 1'b1; frame3.error[ 647] = 1'b0;frame3.data[ 648] = 8'h7C; frame3.valid[ 648] = 1'b1; frame3.error[ 648] = 1'b0;frame3.data[ 649] = 8'h7D; frame3.valid[ 649] = 1'b1; frame3.error[ 649] = 1'b0;frame3.data[ 650] = 8'h7E; frame3.valid[ 650] = 1'b1; frame3.error[ 650] = 1'b0;frame3.data[ 651] = 8'h7F; frame3.valid[ 651] = 1'b1; frame3.error[ 651] = 1'b0;frame3.data[ 652] = 8'h80; frame3.valid[ 652] = 1'b1; frame3.error[ 652] = 1'b0;frame3.data[ 653] = 8'h81; frame3.valid[ 653] = 1'b1; frame3.error[ 653] = 1'b0;
        frame3.data[ 654] = 8'h82; frame3.valid[ 654] = 1'b1; frame3.error[ 654] = 1'b0;frame3.data[ 655] = 8'h83; frame3.valid[ 655] = 1'b1; frame3.error[ 655] = 1'b0;frame3.data[ 656] = 8'h84; frame3.valid[ 656] = 1'b1; frame3.error[ 656] = 1'b0;frame3.data[ 657] = 8'h85; frame3.valid[ 657] = 1'b1; frame3.error[ 657] = 1'b0;frame3.data[ 658] = 8'h86; frame3.valid[ 658] = 1'b1; frame3.error[ 658] = 1'b0;frame3.data[ 659] = 8'h87; frame3.valid[ 659] = 1'b1; frame3.error[ 659] = 1'b0;frame3.data[ 660] = 8'h88; frame3.valid[ 660] = 1'b1; frame3.error[ 660] = 1'b0;frame3.data[ 661] = 8'h89; frame3.valid[ 661] = 1'b1; frame3.error[ 661] = 1'b0;frame3.data[ 662] = 8'h8A; frame3.valid[ 662] = 1'b1; frame3.error[ 662] = 1'b0;frame3.data[ 663] = 8'h8B; frame3.valid[ 663] = 1'b1; frame3.error[ 663] = 1'b0;frame3.data[ 664] = 8'h8C; frame3.valid[ 664] = 1'b1; frame3.error[ 664] = 1'b0;frame3.data[ 665] = 8'h8D; frame3.valid[ 665] = 1'b1; frame3.error[ 665] = 1'b0;frame3.data[ 666] = 8'h8E; frame3.valid[ 666] = 1'b1; frame3.error[ 666] = 1'b0;frame3.data[ 667] = 8'h8F; frame3.valid[ 667] = 1'b1; frame3.error[ 667] = 1'b0;frame3.data[ 668] = 8'h90; frame3.valid[ 668] = 1'b1; frame3.error[ 668] = 1'b0;frame3.data[ 669] = 8'h91; frame3.valid[ 669] = 1'b1; frame3.error[ 669] = 1'b0;
        frame3.data[ 670] = 8'h92; frame3.valid[ 670] = 1'b1; frame3.error[ 670] = 1'b0;frame3.data[ 671] = 8'h93; frame3.valid[ 671] = 1'b1; frame3.error[ 671] = 1'b0;frame3.data[ 672] = 8'h94; frame3.valid[ 672] = 1'b1; frame3.error[ 672] = 1'b0;frame3.data[ 673] = 8'h95; frame3.valid[ 673] = 1'b1; frame3.error[ 673] = 1'b0;frame3.data[ 674] = 8'h96; frame3.valid[ 674] = 1'b1; frame3.error[ 674] = 1'b0;frame3.data[ 675] = 8'h97; frame3.valid[ 675] = 1'b1; frame3.error[ 675] = 1'b0;frame3.data[ 676] = 8'h98; frame3.valid[ 676] = 1'b1; frame3.error[ 676] = 1'b0;frame3.data[ 677] = 8'h99; frame3.valid[ 677] = 1'b1; frame3.error[ 677] = 1'b0;frame3.data[ 678] = 8'h9A; frame3.valid[ 678] = 1'b1; frame3.error[ 678] = 1'b0;frame3.data[ 679] = 8'h9B; frame3.valid[ 679] = 1'b1; frame3.error[ 679] = 1'b0;frame3.data[ 680] = 8'h9C; frame3.valid[ 680] = 1'b1; frame3.error[ 680] = 1'b0;frame3.data[ 681] = 8'h9D; frame3.valid[ 681] = 1'b1; frame3.error[ 681] = 1'b0;frame3.data[ 682] = 8'h9E; frame3.valid[ 682] = 1'b1; frame3.error[ 682] = 1'b0;frame3.data[ 683] = 8'h9F; frame3.valid[ 683] = 1'b1; frame3.error[ 683] = 1'b0;frame3.data[ 684] = 8'hA0; frame3.valid[ 684] = 1'b1; frame3.error[ 684] = 1'b0;frame3.data[ 685] = 8'hA1; frame3.valid[ 685] = 1'b1; frame3.error[ 685] = 1'b0;
        frame3.data[ 686] = 8'hA2; frame3.valid[ 686] = 1'b1; frame3.error[ 686] = 1'b0;frame3.data[ 687] = 8'hA3; frame3.valid[ 687] = 1'b1; frame3.error[ 687] = 1'b0;frame3.data[ 688] = 8'hA4; frame3.valid[ 688] = 1'b1; frame3.error[ 688] = 1'b0;frame3.data[ 689] = 8'hA5; frame3.valid[ 689] = 1'b1; frame3.error[ 689] = 1'b0;frame3.data[ 690] = 8'hA6; frame3.valid[ 690] = 1'b1; frame3.error[ 690] = 1'b0;frame3.data[ 691] = 8'hA7; frame3.valid[ 691] = 1'b1; frame3.error[ 691] = 1'b0;frame3.data[ 692] = 8'hA8; frame3.valid[ 692] = 1'b1; frame3.error[ 692] = 1'b0;frame3.data[ 693] = 8'hA9; frame3.valid[ 693] = 1'b1; frame3.error[ 693] = 1'b0;frame3.data[ 694] = 8'hAA; frame3.valid[ 694] = 1'b1; frame3.error[ 694] = 1'b0;frame3.data[ 695] = 8'hAB; frame3.valid[ 695] = 1'b1; frame3.error[ 695] = 1'b0;frame3.data[ 696] = 8'hAC; frame3.valid[ 696] = 1'b1; frame3.error[ 696] = 1'b0;frame3.data[ 697] = 8'hAD; frame3.valid[ 697] = 1'b1; frame3.error[ 697] = 1'b0;frame3.data[ 698] = 8'hAE; frame3.valid[ 698] = 1'b1; frame3.error[ 698] = 1'b0;frame3.data[ 699] = 8'hAF; frame3.valid[ 699] = 1'b1; frame3.error[ 699] = 1'b0;frame3.data[ 700] = 8'hB0; frame3.valid[ 700] = 1'b1; frame3.error[ 700] = 1'b0;frame3.data[ 701] = 8'hB1; frame3.valid[ 701] = 1'b1; frame3.error[ 701] = 1'b0;
        frame3.data[ 702] = 8'hB2; frame3.valid[ 702] = 1'b1; frame3.error[ 702] = 1'b0;frame3.data[ 703] = 8'hB3; frame3.valid[ 703] = 1'b1; frame3.error[ 703] = 1'b0;frame3.data[ 704] = 8'hB4; frame3.valid[ 704] = 1'b1; frame3.error[ 704] = 1'b0;frame3.data[ 705] = 8'hB5; frame3.valid[ 705] = 1'b1; frame3.error[ 705] = 1'b0;frame3.data[ 706] = 8'hB6; frame3.valid[ 706] = 1'b1; frame3.error[ 706] = 1'b0;frame3.data[ 707] = 8'hB7; frame3.valid[ 707] = 1'b1; frame3.error[ 707] = 1'b0;frame3.data[ 708] = 8'hB8; frame3.valid[ 708] = 1'b1; frame3.error[ 708] = 1'b0;frame3.data[ 709] = 8'hB9; frame3.valid[ 709] = 1'b1; frame3.error[ 709] = 1'b0;frame3.data[ 710] = 8'hBA; frame3.valid[ 710] = 1'b1; frame3.error[ 710] = 1'b0;frame3.data[ 711] = 8'hBB; frame3.valid[ 711] = 1'b1; frame3.error[ 711] = 1'b0;frame3.data[ 712] = 8'hBC; frame3.valid[ 712] = 1'b1; frame3.error[ 712] = 1'b0;frame3.data[ 713] = 8'hBD; frame3.valid[ 713] = 1'b1; frame3.error[ 713] = 1'b0;frame3.data[ 714] = 8'hBE; frame3.valid[ 714] = 1'b1; frame3.error[ 714] = 1'b0;frame3.data[ 715] = 8'hBF; frame3.valid[ 715] = 1'b1; frame3.error[ 715] = 1'b0;frame3.data[ 716] = 8'hC0; frame3.valid[ 716] = 1'b1; frame3.error[ 716] = 1'b0;frame3.data[ 717] = 8'hC1; frame3.valid[ 717] = 1'b1; frame3.error[ 717] = 1'b0;
        frame3.data[ 718] = 8'hC2; frame3.valid[ 718] = 1'b1; frame3.error[ 718] = 1'b0;frame3.data[ 719] = 8'hC3; frame3.valid[ 719] = 1'b1; frame3.error[ 719] = 1'b0;frame3.data[ 720] = 8'hC4; frame3.valid[ 720] = 1'b1; frame3.error[ 720] = 1'b0;frame3.data[ 721] = 8'hC5; frame3.valid[ 721] = 1'b1; frame3.error[ 721] = 1'b0;frame3.data[ 722] = 8'hC6; frame3.valid[ 722] = 1'b1; frame3.error[ 722] = 1'b0;frame3.data[ 723] = 8'hC7; frame3.valid[ 723] = 1'b1; frame3.error[ 723] = 1'b0;frame3.data[ 724] = 8'hC8; frame3.valid[ 724] = 1'b1; frame3.error[ 724] = 1'b0;frame3.data[ 725] = 8'hC9; frame3.valid[ 725] = 1'b1; frame3.error[ 725] = 1'b0;frame3.data[ 726] = 8'hCA; frame3.valid[ 726] = 1'b1; frame3.error[ 726] = 1'b0;frame3.data[ 727] = 8'hCB; frame3.valid[ 727] = 1'b1; frame3.error[ 727] = 1'b0;frame3.data[ 728] = 8'hCC; frame3.valid[ 728] = 1'b1; frame3.error[ 728] = 1'b0;frame3.data[ 729] = 8'hCD; frame3.valid[ 729] = 1'b1; frame3.error[ 729] = 1'b0;frame3.data[ 730] = 8'hCE; frame3.valid[ 730] = 1'b1; frame3.error[ 730] = 1'b0;frame3.data[ 731] = 8'hCF; frame3.valid[ 731] = 1'b1; frame3.error[ 731] = 1'b0;frame3.data[ 732] = 8'hD0; frame3.valid[ 732] = 1'b1; frame3.error[ 732] = 1'b0;frame3.data[ 733] = 8'hD1; frame3.valid[ 733] = 1'b1; frame3.error[ 733] = 1'b0;
        frame3.data[ 734] = 8'hD2; frame3.valid[ 734] = 1'b1; frame3.error[ 734] = 1'b0;frame3.data[ 735] = 8'hD3; frame3.valid[ 735] = 1'b1; frame3.error[ 735] = 1'b0;frame3.data[ 736] = 8'hD4; frame3.valid[ 736] = 1'b1; frame3.error[ 736] = 1'b0;frame3.data[ 737] = 8'hD5; frame3.valid[ 737] = 1'b1; frame3.error[ 737] = 1'b0;frame3.data[ 738] = 8'hD6; frame3.valid[ 738] = 1'b1; frame3.error[ 738] = 1'b0;frame3.data[ 739] = 8'hD7; frame3.valid[ 739] = 1'b1; frame3.error[ 739] = 1'b0;frame3.data[ 740] = 8'hD8; frame3.valid[ 740] = 1'b1; frame3.error[ 740] = 1'b0;frame3.data[ 741] = 8'hD9; frame3.valid[ 741] = 1'b1; frame3.error[ 741] = 1'b0;frame3.data[ 742] = 8'hDA; frame3.valid[ 742] = 1'b1; frame3.error[ 742] = 1'b0;frame3.data[ 743] = 8'hDB; frame3.valid[ 743] = 1'b1; frame3.error[ 743] = 1'b0;frame3.data[ 744] = 8'hDC; frame3.valid[ 744] = 1'b1; frame3.error[ 744] = 1'b0;frame3.data[ 745] = 8'hDD; frame3.valid[ 745] = 1'b1; frame3.error[ 745] = 1'b0;frame3.data[ 746] = 8'hDE; frame3.valid[ 746] = 1'b1; frame3.error[ 746] = 1'b0;frame3.data[ 747] = 8'hDF; frame3.valid[ 747] = 1'b1; frame3.error[ 747] = 1'b0;frame3.data[ 748] = 8'hE0; frame3.valid[ 748] = 1'b1; frame3.error[ 748] = 1'b0;frame3.data[ 749] = 8'hE1; frame3.valid[ 749] = 1'b1; frame3.error[ 749] = 1'b0;
        frame3.data[ 750] = 8'hE2; frame3.valid[ 750] = 1'b1; frame3.error[ 750] = 1'b0;frame3.data[ 751] = 8'hE3; frame3.valid[ 751] = 1'b1; frame3.error[ 751] = 1'b0;frame3.data[ 752] = 8'hE4; frame3.valid[ 752] = 1'b1; frame3.error[ 752] = 1'b0;frame3.data[ 753] = 8'hE5; frame3.valid[ 753] = 1'b1; frame3.error[ 753] = 1'b0;frame3.data[ 754] = 8'hE6; frame3.valid[ 754] = 1'b1; frame3.error[ 754] = 1'b0;frame3.data[ 755] = 8'hE7; frame3.valid[ 755] = 1'b1; frame3.error[ 755] = 1'b0;frame3.data[ 756] = 8'hE8; frame3.valid[ 756] = 1'b1; frame3.error[ 756] = 1'b0;frame3.data[ 757] = 8'hE9; frame3.valid[ 757] = 1'b1; frame3.error[ 757] = 1'b0;frame3.data[ 758] = 8'hEA; frame3.valid[ 758] = 1'b1; frame3.error[ 758] = 1'b0;frame3.data[ 759] = 8'hEB; frame3.valid[ 759] = 1'b1; frame3.error[ 759] = 1'b0;frame3.data[ 760] = 8'hEC; frame3.valid[ 760] = 1'b1; frame3.error[ 760] = 1'b0;frame3.data[ 761] = 8'hED; frame3.valid[ 761] = 1'b1; frame3.error[ 761] = 1'b0;frame3.data[ 762] = 8'hEE; frame3.valid[ 762] = 1'b1; frame3.error[ 762] = 1'b0;frame3.data[ 763] = 8'hEF; frame3.valid[ 763] = 1'b1; frame3.error[ 763] = 1'b0;frame3.data[ 764] = 8'hF0; frame3.valid[ 764] = 1'b1; frame3.error[ 764] = 1'b0;frame3.data[ 765] = 8'hF1; frame3.valid[ 765] = 1'b1; frame3.error[ 765] = 1'b0;
        frame3.data[ 766] = 8'hF2; frame3.valid[ 766] = 1'b1; frame3.error[ 766] = 1'b0;frame3.data[ 767] = 8'hF3; frame3.valid[ 767] = 1'b1; frame3.error[ 767] = 1'b0;frame3.data[ 768] = 8'hF4; frame3.valid[ 768] = 1'b1; frame3.error[ 768] = 1'b0;frame3.data[ 769] = 8'hF5; frame3.valid[ 769] = 1'b1; frame3.error[ 769] = 1'b0;frame3.data[ 770] = 8'hF6; frame3.valid[ 770] = 1'b1; frame3.error[ 770] = 1'b0;frame3.data[ 771] = 8'hF7; frame3.valid[ 771] = 1'b1; frame3.error[ 771] = 1'b0;frame3.data[ 772] = 8'hF8; frame3.valid[ 772] = 1'b1; frame3.error[ 772] = 1'b0;frame3.data[ 773] = 8'hF9; frame3.valid[ 773] = 1'b1; frame3.error[ 773] = 1'b0;frame3.data[ 774] = 8'hFA; frame3.valid[ 774] = 1'b1; frame3.error[ 774] = 1'b0;frame3.data[ 775] = 8'hFB; frame3.valid[ 775] = 1'b1; frame3.error[ 775] = 1'b0;frame3.data[ 776] = 8'hFC; frame3.valid[ 776] = 1'b1; frame3.error[ 776] = 1'b0;frame3.data[ 777] = 8'hFD; frame3.valid[ 777] = 1'b1; frame3.error[ 777] = 1'b0;frame3.data[ 778] = 8'hFE; frame3.valid[ 778] = 1'b1; frame3.error[ 778] = 1'b0;frame3.data[ 779] = 8'h00; frame3.valid[ 779] = 1'b1; frame3.error[ 779] = 1'b0;frame3.data[ 780] = 8'h01; frame3.valid[ 780] = 1'b1; frame3.error[ 780] = 1'b0;frame3.data[ 781] = 8'h02; frame3.valid[ 781] = 1'b1; frame3.error[ 781] = 1'b0;
        frame3.data[ 782] = 8'h03; frame3.valid[ 782] = 1'b1; frame3.error[ 782] = 1'b0;frame3.data[ 783] = 8'h04; frame3.valid[ 783] = 1'b1; frame3.error[ 783] = 1'b0;frame3.data[ 784] = 8'h05; frame3.valid[ 784] = 1'b1; frame3.error[ 784] = 1'b0;frame3.data[ 785] = 8'h06; frame3.valid[ 785] = 1'b1; frame3.error[ 785] = 1'b0;frame3.data[ 786] = 8'h07; frame3.valid[ 786] = 1'b1; frame3.error[ 786] = 1'b0;frame3.data[ 787] = 8'h08; frame3.valid[ 787] = 1'b1; frame3.error[ 787] = 1'b0;frame3.data[ 788] = 8'h09; frame3.valid[ 788] = 1'b1; frame3.error[ 788] = 1'b0;frame3.data[ 789] = 8'h0A; frame3.valid[ 789] = 1'b1; frame3.error[ 789] = 1'b0;frame3.data[ 790] = 8'h0B; frame3.valid[ 790] = 1'b1; frame3.error[ 790] = 1'b0;frame3.data[ 791] = 8'h0C; frame3.valid[ 791] = 1'b1; frame3.error[ 791] = 1'b0;frame3.data[ 792] = 8'h0D; frame3.valid[ 792] = 1'b1; frame3.error[ 792] = 1'b0;frame3.data[ 793] = 8'h0E; frame3.valid[ 793] = 1'b1; frame3.error[ 793] = 1'b0;frame3.data[ 794] = 8'h0F; frame3.valid[ 794] = 1'b1; frame3.error[ 794] = 1'b0;frame3.data[ 795] = 8'h10; frame3.valid[ 795] = 1'b1; frame3.error[ 795] = 1'b0;frame3.data[ 796] = 8'h11; frame3.valid[ 796] = 1'b1; frame3.error[ 796] = 1'b0;frame3.data[ 797] = 8'h12; frame3.valid[ 797] = 1'b1; frame3.error[ 797] = 1'b0;
        frame3.data[ 798] = 8'h13; frame3.valid[ 798] = 1'b1; frame3.error[ 798] = 1'b0;frame3.data[ 799] = 8'h14; frame3.valid[ 799] = 1'b1; frame3.error[ 799] = 1'b0;frame3.data[ 800] = 8'h15; frame3.valid[ 800] = 1'b1; frame3.error[ 800] = 1'b0;frame3.data[ 801] = 8'h16; frame3.valid[ 801] = 1'b1; frame3.error[ 801] = 1'b0;frame3.data[ 802] = 8'h17; frame3.valid[ 802] = 1'b1; frame3.error[ 802] = 1'b0;frame3.data[ 803] = 8'h18; frame3.valid[ 803] = 1'b1; frame3.error[ 803] = 1'b0;frame3.data[ 804] = 8'h19; frame3.valid[ 804] = 1'b1; frame3.error[ 804] = 1'b0;frame3.data[ 805] = 8'h1A; frame3.valid[ 805] = 1'b1; frame3.error[ 805] = 1'b0;frame3.data[ 806] = 8'h1B; frame3.valid[ 806] = 1'b1; frame3.error[ 806] = 1'b0;frame3.data[ 807] = 8'h1C; frame3.valid[ 807] = 1'b1; frame3.error[ 807] = 1'b0;frame3.data[ 808] = 8'h1D; frame3.valid[ 808] = 1'b1; frame3.error[ 808] = 1'b0;frame3.data[ 809] = 8'h1E; frame3.valid[ 809] = 1'b1; frame3.error[ 809] = 1'b0;frame3.data[ 810] = 8'h1F; frame3.valid[ 810] = 1'b1; frame3.error[ 810] = 1'b0;frame3.data[ 811] = 8'h20; frame3.valid[ 811] = 1'b1; frame3.error[ 811] = 1'b0;frame3.data[ 812] = 8'h21; frame3.valid[ 812] = 1'b1; frame3.error[ 812] = 1'b0;frame3.data[ 813] = 8'h22; frame3.valid[ 813] = 1'b1; frame3.error[ 813] = 1'b0;
        frame3.data[ 814] = 8'h23; frame3.valid[ 814] = 1'b1; frame3.error[ 814] = 1'b0;frame3.data[ 815] = 8'h24; frame3.valid[ 815] = 1'b1; frame3.error[ 815] = 1'b0;frame3.data[ 816] = 8'h25; frame3.valid[ 816] = 1'b1; frame3.error[ 816] = 1'b0;frame3.data[ 817] = 8'h26; frame3.valid[ 817] = 1'b1; frame3.error[ 817] = 1'b0;frame3.data[ 818] = 8'h27; frame3.valid[ 818] = 1'b1; frame3.error[ 818] = 1'b0;frame3.data[ 819] = 8'h28; frame3.valid[ 819] = 1'b1; frame3.error[ 819] = 1'b0;frame3.data[ 820] = 8'h29; frame3.valid[ 820] = 1'b1; frame3.error[ 820] = 1'b0;frame3.data[ 821] = 8'h2A; frame3.valid[ 821] = 1'b1; frame3.error[ 821] = 1'b0;frame3.data[ 822] = 8'h2B; frame3.valid[ 822] = 1'b1; frame3.error[ 822] = 1'b0;frame3.data[ 823] = 8'h2C; frame3.valid[ 823] = 1'b1; frame3.error[ 823] = 1'b0;frame3.data[ 824] = 8'h2D; frame3.valid[ 824] = 1'b1; frame3.error[ 824] = 1'b0;frame3.data[ 825] = 8'h2E; frame3.valid[ 825] = 1'b1; frame3.error[ 825] = 1'b0;frame3.data[ 826] = 8'h2F; frame3.valid[ 826] = 1'b1; frame3.error[ 826] = 1'b0;frame3.data[ 827] = 8'h30; frame3.valid[ 827] = 1'b1; frame3.error[ 827] = 1'b0;frame3.data[ 828] = 8'h31; frame3.valid[ 828] = 1'b1; frame3.error[ 828] = 1'b0;frame3.data[ 829] = 8'h32; frame3.valid[ 829] = 1'b1; frame3.error[ 829] = 1'b0;
        frame3.data[ 830] = 8'h33; frame3.valid[ 830] = 1'b1; frame3.error[ 830] = 1'b0;frame3.data[ 831] = 8'h34; frame3.valid[ 831] = 1'b1; frame3.error[ 831] = 1'b0;frame3.data[ 832] = 8'h35; frame3.valid[ 832] = 1'b1; frame3.error[ 832] = 1'b0;frame3.data[ 833] = 8'h36; frame3.valid[ 833] = 1'b1; frame3.error[ 833] = 1'b0;frame3.data[ 834] = 8'h37; frame3.valid[ 834] = 1'b1; frame3.error[ 834] = 1'b0;frame3.data[ 835] = 8'h38; frame3.valid[ 835] = 1'b1; frame3.error[ 835] = 1'b0;frame3.data[ 836] = 8'h39; frame3.valid[ 836] = 1'b1; frame3.error[ 836] = 1'b0;frame3.data[ 837] = 8'h3A; frame3.valid[ 837] = 1'b1; frame3.error[ 837] = 1'b0;frame3.data[ 838] = 8'h3B; frame3.valid[ 838] = 1'b1; frame3.error[ 838] = 1'b0;frame3.data[ 839] = 8'h3C; frame3.valid[ 839] = 1'b1; frame3.error[ 839] = 1'b0;frame3.data[ 840] = 8'h3D; frame3.valid[ 840] = 1'b1; frame3.error[ 840] = 1'b0;frame3.data[ 841] = 8'h3E; frame3.valid[ 841] = 1'b1; frame3.error[ 841] = 1'b0;frame3.data[ 842] = 8'h3F; frame3.valid[ 842] = 1'b1; frame3.error[ 842] = 1'b0;frame3.data[ 843] = 8'h40; frame3.valid[ 843] = 1'b1; frame3.error[ 843] = 1'b0;frame3.data[ 844] = 8'h41; frame3.valid[ 844] = 1'b1; frame3.error[ 844] = 1'b0;frame3.data[ 845] = 8'h42; frame3.valid[ 845] = 1'b1; frame3.error[ 845] = 1'b0;
        frame3.data[ 846] = 8'h43; frame3.valid[ 846] = 1'b1; frame3.error[ 846] = 1'b0;frame3.data[ 847] = 8'h44; frame3.valid[ 847] = 1'b1; frame3.error[ 847] = 1'b0;frame3.data[ 848] = 8'h45; frame3.valid[ 848] = 1'b1; frame3.error[ 848] = 1'b0;frame3.data[ 849] = 8'h46; frame3.valid[ 849] = 1'b1; frame3.error[ 849] = 1'b0;frame3.data[ 850] = 8'h47; frame3.valid[ 850] = 1'b1; frame3.error[ 850] = 1'b0;frame3.data[ 851] = 8'h48; frame3.valid[ 851] = 1'b1; frame3.error[ 851] = 1'b0;frame3.data[ 852] = 8'h49; frame3.valid[ 852] = 1'b1; frame3.error[ 852] = 1'b0;frame3.data[ 853] = 8'h4A; frame3.valid[ 853] = 1'b1; frame3.error[ 853] = 1'b0;frame3.data[ 854] = 8'h4B; frame3.valid[ 854] = 1'b1; frame3.error[ 854] = 1'b0;frame3.data[ 855] = 8'h4C; frame3.valid[ 855] = 1'b1; frame3.error[ 855] = 1'b0;frame3.data[ 856] = 8'h4D; frame3.valid[ 856] = 1'b1; frame3.error[ 856] = 1'b0;frame3.data[ 857] = 8'h4E; frame3.valid[ 857] = 1'b1; frame3.error[ 857] = 1'b0;frame3.data[ 858] = 8'h4F; frame3.valid[ 858] = 1'b1; frame3.error[ 858] = 1'b0;frame3.data[ 859] = 8'h50; frame3.valid[ 859] = 1'b1; frame3.error[ 859] = 1'b0;frame3.data[ 860] = 8'h51; frame3.valid[ 860] = 1'b1; frame3.error[ 860] = 1'b0;frame3.data[ 861] = 8'h52; frame3.valid[ 861] = 1'b1; frame3.error[ 861] = 1'b0;
        frame3.data[ 862] = 8'h53; frame3.valid[ 862] = 1'b1; frame3.error[ 862] = 1'b0;frame3.data[ 863] = 8'h54; frame3.valid[ 863] = 1'b1; frame3.error[ 863] = 1'b0;frame3.data[ 864] = 8'h55; frame3.valid[ 864] = 1'b1; frame3.error[ 864] = 1'b0;frame3.data[ 865] = 8'h56; frame3.valid[ 865] = 1'b1; frame3.error[ 865] = 1'b0;frame3.data[ 866] = 8'h57; frame3.valid[ 866] = 1'b1; frame3.error[ 866] = 1'b0;frame3.data[ 867] = 8'h58; frame3.valid[ 867] = 1'b1; frame3.error[ 867] = 1'b0;frame3.data[ 868] = 8'h59; frame3.valid[ 868] = 1'b1; frame3.error[ 868] = 1'b0;frame3.data[ 869] = 8'h5A; frame3.valid[ 869] = 1'b1; frame3.error[ 869] = 1'b0;frame3.data[ 870] = 8'h5B; frame3.valid[ 870] = 1'b1; frame3.error[ 870] = 1'b0;frame3.data[ 871] = 8'h5C; frame3.valid[ 871] = 1'b1; frame3.error[ 871] = 1'b0;frame3.data[ 872] = 8'h5D; frame3.valid[ 872] = 1'b1; frame3.error[ 872] = 1'b0;frame3.data[ 873] = 8'h5E; frame3.valid[ 873] = 1'b1; frame3.error[ 873] = 1'b0;frame3.data[ 874] = 8'h5F; frame3.valid[ 874] = 1'b1; frame3.error[ 874] = 1'b0;frame3.data[ 875] = 8'h60; frame3.valid[ 875] = 1'b1; frame3.error[ 875] = 1'b0;frame3.data[ 876] = 8'h61; frame3.valid[ 876] = 1'b1; frame3.error[ 876] = 1'b0;frame3.data[ 877] = 8'h62; frame3.valid[ 877] = 1'b1; frame3.error[ 877] = 1'b0;
        frame3.data[ 878] = 8'h63; frame3.valid[ 878] = 1'b1; frame3.error[ 878] = 1'b0;frame3.data[ 879] = 8'h64; frame3.valid[ 879] = 1'b1; frame3.error[ 879] = 1'b0;frame3.data[ 880] = 8'h65; frame3.valid[ 880] = 1'b1; frame3.error[ 880] = 1'b0;frame3.data[ 881] = 8'h66; frame3.valid[ 881] = 1'b1; frame3.error[ 881] = 1'b0;frame3.data[ 882] = 8'h67; frame3.valid[ 882] = 1'b1; frame3.error[ 882] = 1'b0;frame3.data[ 883] = 8'h68; frame3.valid[ 883] = 1'b1; frame3.error[ 883] = 1'b0;frame3.data[ 884] = 8'h69; frame3.valid[ 884] = 1'b1; frame3.error[ 884] = 1'b0;frame3.data[ 885] = 8'h6A; frame3.valid[ 885] = 1'b1; frame3.error[ 885] = 1'b0;frame3.data[ 886] = 8'h6B; frame3.valid[ 886] = 1'b1; frame3.error[ 886] = 1'b0;frame3.data[ 887] = 8'h6C; frame3.valid[ 887] = 1'b1; frame3.error[ 887] = 1'b0;frame3.data[ 888] = 8'h6D; frame3.valid[ 888] = 1'b1; frame3.error[ 888] = 1'b0;frame3.data[ 889] = 8'h6E; frame3.valid[ 889] = 1'b1; frame3.error[ 889] = 1'b0;frame3.data[ 890] = 8'h6F; frame3.valid[ 890] = 1'b1; frame3.error[ 890] = 1'b0;frame3.data[ 891] = 8'h70; frame3.valid[ 891] = 1'b1; frame3.error[ 891] = 1'b0;frame3.data[ 892] = 8'h71; frame3.valid[ 892] = 1'b1; frame3.error[ 892] = 1'b0;frame3.data[ 893] = 8'h72; frame3.valid[ 893] = 1'b1; frame3.error[ 893] = 1'b0;
        frame3.data[ 894] = 8'h73; frame3.valid[ 894] = 1'b1; frame3.error[ 894] = 1'b0;frame3.data[ 895] = 8'h74; frame3.valid[ 895] = 1'b1; frame3.error[ 895] = 1'b0;frame3.data[ 896] = 8'h75; frame3.valid[ 896] = 1'b1; frame3.error[ 896] = 1'b0;frame3.data[ 897] = 8'h76; frame3.valid[ 897] = 1'b1; frame3.error[ 897] = 1'b0;frame3.data[ 898] = 8'h77; frame3.valid[ 898] = 1'b1; frame3.error[ 898] = 1'b0;frame3.data[ 899] = 8'h78; frame3.valid[ 899] = 1'b1; frame3.error[ 899] = 1'b0;frame3.data[ 900] = 8'h79; frame3.valid[ 900] = 1'b1; frame3.error[ 900] = 1'b0;frame3.data[ 901] = 8'h7A; frame3.valid[ 901] = 1'b1; frame3.error[ 901] = 1'b0;frame3.data[ 902] = 8'h7B; frame3.valid[ 902] = 1'b1; frame3.error[ 902] = 1'b0;frame3.data[ 903] = 8'h7C; frame3.valid[ 903] = 1'b1; frame3.error[ 903] = 1'b0;frame3.data[ 904] = 8'h7D; frame3.valid[ 904] = 1'b1; frame3.error[ 904] = 1'b0;frame3.data[ 905] = 8'h7E; frame3.valid[ 905] = 1'b1; frame3.error[ 905] = 1'b0;frame3.data[ 906] = 8'h7F; frame3.valid[ 906] = 1'b1; frame3.error[ 906] = 1'b0;frame3.data[ 907] = 8'h80; frame3.valid[ 907] = 1'b1; frame3.error[ 907] = 1'b0;frame3.data[ 908] = 8'h81; frame3.valid[ 908] = 1'b1; frame3.error[ 908] = 1'b0;frame3.data[ 909] = 8'h82; frame3.valid[ 909] = 1'b1; frame3.error[ 909] = 1'b0;
        frame3.data[ 910] = 8'h83; frame3.valid[ 910] = 1'b1; frame3.error[ 910] = 1'b0;frame3.data[ 911] = 8'h84; frame3.valid[ 911] = 1'b1; frame3.error[ 911] = 1'b0;frame3.data[ 912] = 8'h85; frame3.valid[ 912] = 1'b1; frame3.error[ 912] = 1'b0;frame3.data[ 913] = 8'h86; frame3.valid[ 913] = 1'b1; frame3.error[ 913] = 1'b0;frame3.data[ 914] = 8'h87; frame3.valid[ 914] = 1'b1; frame3.error[ 914] = 1'b0;frame3.data[ 915] = 8'h88; frame3.valid[ 915] = 1'b1; frame3.error[ 915] = 1'b0;frame3.data[ 916] = 8'h89; frame3.valid[ 916] = 1'b1; frame3.error[ 916] = 1'b0;frame3.data[ 917] = 8'h8A; frame3.valid[ 917] = 1'b1; frame3.error[ 917] = 1'b0;frame3.data[ 918] = 8'h8B; frame3.valid[ 918] = 1'b1; frame3.error[ 918] = 1'b0;frame3.data[ 919] = 8'h8C; frame3.valid[ 919] = 1'b1; frame3.error[ 919] = 1'b0;frame3.data[ 920] = 8'h8D; frame3.valid[ 920] = 1'b1; frame3.error[ 920] = 1'b0;frame3.data[ 921] = 8'h8E; frame3.valid[ 921] = 1'b1; frame3.error[ 921] = 1'b0;frame3.data[ 922] = 8'h8F; frame3.valid[ 922] = 1'b1; frame3.error[ 922] = 1'b0;frame3.data[ 923] = 8'h90; frame3.valid[ 923] = 1'b1; frame3.error[ 923] = 1'b0;frame3.data[ 924] = 8'h91; frame3.valid[ 924] = 1'b1; frame3.error[ 924] = 1'b0;frame3.data[ 925] = 8'h92; frame3.valid[ 925] = 1'b1; frame3.error[ 925] = 1'b0;
        frame3.data[ 926] = 8'h93; frame3.valid[ 926] = 1'b1; frame3.error[ 926] = 1'b0;frame3.data[ 927] = 8'h94; frame3.valid[ 927] = 1'b1; frame3.error[ 927] = 1'b0;frame3.data[ 928] = 8'h95; frame3.valid[ 928] = 1'b1; frame3.error[ 928] = 1'b0;frame3.data[ 929] = 8'h96; frame3.valid[ 929] = 1'b1; frame3.error[ 929] = 1'b0;frame3.data[ 930] = 8'h97; frame3.valid[ 930] = 1'b1; frame3.error[ 930] = 1'b0;frame3.data[ 931] = 8'h98; frame3.valid[ 931] = 1'b1; frame3.error[ 931] = 1'b0;frame3.data[ 932] = 8'h99; frame3.valid[ 932] = 1'b1; frame3.error[ 932] = 1'b0;frame3.data[ 933] = 8'h9A; frame3.valid[ 933] = 1'b1; frame3.error[ 933] = 1'b0;frame3.data[ 934] = 8'h9B; frame3.valid[ 934] = 1'b1; frame3.error[ 934] = 1'b0;frame3.data[ 935] = 8'h9C; frame3.valid[ 935] = 1'b1; frame3.error[ 935] = 1'b0;frame3.data[ 936] = 8'h9D; frame3.valid[ 936] = 1'b1; frame3.error[ 936] = 1'b0;frame3.data[ 937] = 8'h9E; frame3.valid[ 937] = 1'b1; frame3.error[ 937] = 1'b0;frame3.data[ 938] = 8'h9F; frame3.valid[ 938] = 1'b1; frame3.error[ 938] = 1'b0;frame3.data[ 939] = 8'hA0; frame3.valid[ 939] = 1'b1; frame3.error[ 939] = 1'b0;frame3.data[ 940] = 8'hA1; frame3.valid[ 940] = 1'b1; frame3.error[ 940] = 1'b0;frame3.data[ 941] = 8'hA2; frame3.valid[ 941] = 1'b1; frame3.error[ 941] = 1'b0;
        frame3.data[ 942] = 8'hA3; frame3.valid[ 942] = 1'b1; frame3.error[ 942] = 1'b0;frame3.data[ 943] = 8'hA4; frame3.valid[ 943] = 1'b1; frame3.error[ 943] = 1'b0;frame3.data[ 944] = 8'hA5; frame3.valid[ 944] = 1'b1; frame3.error[ 944] = 1'b0;frame3.data[ 945] = 8'hA6; frame3.valid[ 945] = 1'b1; frame3.error[ 945] = 1'b0;frame3.data[ 946] = 8'hA7; frame3.valid[ 946] = 1'b1; frame3.error[ 946] = 1'b0;frame3.data[ 947] = 8'hA8; frame3.valid[ 947] = 1'b1; frame3.error[ 947] = 1'b0;frame3.data[ 948] = 8'hA9; frame3.valid[ 948] = 1'b1; frame3.error[ 948] = 1'b0;frame3.data[ 949] = 8'hAA; frame3.valid[ 949] = 1'b1; frame3.error[ 949] = 1'b0;frame3.data[ 950] = 8'hAB; frame3.valid[ 950] = 1'b1; frame3.error[ 950] = 1'b0;frame3.data[ 951] = 8'hAC; frame3.valid[ 951] = 1'b1; frame3.error[ 951] = 1'b0;frame3.data[ 952] = 8'hAD; frame3.valid[ 952] = 1'b1; frame3.error[ 952] = 1'b0;frame3.data[ 953] = 8'hAE; frame3.valid[ 953] = 1'b1; frame3.error[ 953] = 1'b0;frame3.data[ 954] = 8'hAF; frame3.valid[ 954] = 1'b1; frame3.error[ 954] = 1'b0;frame3.data[ 955] = 8'hB0; frame3.valid[ 955] = 1'b1; frame3.error[ 955] = 1'b0;frame3.data[ 956] = 8'hB1; frame3.valid[ 956] = 1'b1; frame3.error[ 956] = 1'b0;frame3.data[ 957] = 8'hB2; frame3.valid[ 957] = 1'b1; frame3.error[ 957] = 1'b0;
        frame3.data[ 958] = 8'hB3; frame3.valid[ 958] = 1'b1; frame3.error[ 958] = 1'b0;frame3.data[ 959] = 8'hB4; frame3.valid[ 959] = 1'b1; frame3.error[ 959] = 1'b0;frame3.data[ 960] = 8'hB5; frame3.valid[ 960] = 1'b1; frame3.error[ 960] = 1'b0;frame3.data[ 961] = 8'hB6; frame3.valid[ 961] = 1'b1; frame3.error[ 961] = 1'b0;frame3.data[ 962] = 8'hB7; frame3.valid[ 962] = 1'b1; frame3.error[ 962] = 1'b0;frame3.data[ 963] = 8'hB8; frame3.valid[ 963] = 1'b1; frame3.error[ 963] = 1'b0;frame3.data[ 964] = 8'hB9; frame3.valid[ 964] = 1'b1; frame3.error[ 964] = 1'b0;frame3.data[ 965] = 8'hBA; frame3.valid[ 965] = 1'b1; frame3.error[ 965] = 1'b0;frame3.data[ 966] = 8'hBB; frame3.valid[ 966] = 1'b1; frame3.error[ 966] = 1'b0;frame3.data[ 967] = 8'hBC; frame3.valid[ 967] = 1'b1; frame3.error[ 967] = 1'b0;frame3.data[ 968] = 8'hBD; frame3.valid[ 968] = 1'b1; frame3.error[ 968] = 1'b0;frame3.data[ 969] = 8'hBE; frame3.valid[ 969] = 1'b1; frame3.error[ 969] = 1'b0;frame3.data[ 970] = 8'hBF; frame3.valid[ 970] = 1'b1; frame3.error[ 970] = 1'b0;frame3.data[ 971] = 8'hC0; frame3.valid[ 971] = 1'b1; frame3.error[ 971] = 1'b0;frame3.data[ 972] = 8'hC1; frame3.valid[ 972] = 1'b1; frame3.error[ 972] = 1'b0;frame3.data[ 973] = 8'hC2; frame3.valid[ 973] = 1'b1; frame3.error[ 973] = 1'b0;
        frame3.data[ 974] = 8'hC3; frame3.valid[ 974] = 1'b1; frame3.error[ 974] = 1'b0;frame3.data[ 975] = 8'hC4; frame3.valid[ 975] = 1'b1; frame3.error[ 975] = 1'b0;frame3.data[ 976] = 8'hC5; frame3.valid[ 976] = 1'b1; frame3.error[ 976] = 1'b0;frame3.data[ 977] = 8'hC6; frame3.valid[ 977] = 1'b1; frame3.error[ 977] = 1'b0;frame3.data[ 978] = 8'hC7; frame3.valid[ 978] = 1'b1; frame3.error[ 978] = 1'b0;frame3.data[ 979] = 8'hC8; frame3.valid[ 979] = 1'b1; frame3.error[ 979] = 1'b0;frame3.data[ 980] = 8'hC9; frame3.valid[ 980] = 1'b1; frame3.error[ 980] = 1'b0;frame3.data[ 981] = 8'hCA; frame3.valid[ 981] = 1'b1; frame3.error[ 981] = 1'b0;frame3.data[ 982] = 8'hCB; frame3.valid[ 982] = 1'b1; frame3.error[ 982] = 1'b0;frame3.data[ 983] = 8'hCC; frame3.valid[ 983] = 1'b1; frame3.error[ 983] = 1'b0;frame3.data[ 984] = 8'hCD; frame3.valid[ 984] = 1'b1; frame3.error[ 984] = 1'b0;frame3.data[ 985] = 8'hCE; frame3.valid[ 985] = 1'b1; frame3.error[ 985] = 1'b0;frame3.data[ 986] = 8'hCF; frame3.valid[ 986] = 1'b1; frame3.error[ 986] = 1'b0;frame3.data[ 987] = 8'hD0; frame3.valid[ 987] = 1'b1; frame3.error[ 987] = 1'b0;frame3.data[ 988] = 8'hD1; frame3.valid[ 988] = 1'b1; frame3.error[ 988] = 1'b0;frame3.data[ 989] = 8'hD2; frame3.valid[ 989] = 1'b1; frame3.error[ 989] = 1'b0;
        frame3.data[ 990] = 8'hD3; frame3.valid[ 990] = 1'b1; frame3.error[ 990] = 1'b0;frame3.data[ 991] = 8'hD4; frame3.valid[ 991] = 1'b1; frame3.error[ 991] = 1'b0;frame3.data[ 992] = 8'hD5; frame3.valid[ 992] = 1'b1; frame3.error[ 992] = 1'b0;frame3.data[ 993] = 8'hD6; frame3.valid[ 993] = 1'b1; frame3.error[ 993] = 1'b0;frame3.data[ 994] = 8'hD7; frame3.valid[ 994] = 1'b1; frame3.error[ 994] = 1'b0;frame3.data[ 995] = 8'hD8; frame3.valid[ 995] = 1'b1; frame3.error[ 995] = 1'b0;frame3.data[ 996] = 8'hD9; frame3.valid[ 996] = 1'b1; frame3.error[ 996] = 1'b0;frame3.data[ 997] = 8'hDA; frame3.valid[ 997] = 1'b1; frame3.error[ 997] = 1'b0;frame3.data[ 998] = 8'hDB; frame3.valid[ 998] = 1'b1; frame3.error[ 998] = 1'b0;frame3.data[ 999] = 8'hDC; frame3.valid[ 999] = 1'b1; frame3.error[ 999] = 1'b0;frame3.data[1000] = 8'hDD; frame3.valid[1000] = 1'b1; frame3.error[1000] = 1'b0;frame3.data[1001] = 8'hDE; frame3.valid[1001] = 1'b1; frame3.error[1001] = 1'b0;frame3.data[1002] = 8'hDF; frame3.valid[1002] = 1'b1; frame3.error[1002] = 1'b0;frame3.data[1003] = 8'hE0; frame3.valid[1003] = 1'b1; frame3.error[1003] = 1'b0;frame3.data[1004] = 8'hE1; frame3.valid[1004] = 1'b1; frame3.error[1004] = 1'b0;frame3.data[1005] = 8'hE2; frame3.valid[1005] = 1'b1; frame3.error[1005] = 1'b0;
        frame3.data[1006] = 8'hE3; frame3.valid[1006] = 1'b1; frame3.error[1006] = 1'b0;frame3.data[1007] = 8'hE4; frame3.valid[1007] = 1'b1; frame3.error[1007] = 1'b0;frame3.data[1008] = 8'hE5; frame3.valid[1008] = 1'b1; frame3.error[1008] = 1'b0;frame3.data[1009] = 8'hE6; frame3.valid[1009] = 1'b1; frame3.error[1009] = 1'b0;frame3.data[1010] = 8'hE7; frame3.valid[1010] = 1'b1; frame3.error[1010] = 1'b0;frame3.data[1011] = 8'hE8; frame3.valid[1011] = 1'b1; frame3.error[1011] = 1'b0;frame3.data[1012] = 8'hE9; frame3.valid[1012] = 1'b1; frame3.error[1012] = 1'b0;frame3.data[1013] = 8'hEA; frame3.valid[1013] = 1'b1; frame3.error[1013] = 1'b0;frame3.data[1014] = 8'hEB; frame3.valid[1014] = 1'b1; frame3.error[1014] = 1'b0;frame3.data[1015] = 8'hEC; frame3.valid[1015] = 1'b1; frame3.error[1015] = 1'b0;frame3.data[1016] = 8'hED; frame3.valid[1016] = 1'b1; frame3.error[1016] = 1'b0;frame3.data[1017] = 8'hEE; frame3.valid[1017] = 1'b1; frame3.error[1017] = 1'b0;frame3.data[1018] = 8'hEF; frame3.valid[1018] = 1'b1; frame3.error[1018] = 1'b0;frame3.data[1019] = 8'hF0; frame3.valid[1019] = 1'b1; frame3.error[1019] = 1'b0;frame3.data[1020] = 8'hF1; frame3.valid[1020] = 1'b1; frame3.error[1020] = 1'b0;frame3.data[1021] = 8'hF2; frame3.valid[1021] = 1'b1; frame3.error[1021] = 1'b0;
        frame3.data[1022] = 8'hF3; frame3.valid[1022] = 1'b1; frame3.error[1022] = 1'b0;frame3.data[1023] = 8'hF4; frame3.valid[1023] = 1'b1; frame3.error[1023] = 1'b0;frame3.data[1024] = 8'hF5; frame3.valid[1024] = 1'b1; frame3.error[1024] = 1'b0;frame3.data[1025] = 8'hF6; frame3.valid[1025] = 1'b1; frame3.error[1025] = 1'b0;frame3.data[1026] = 8'hF7; frame3.valid[1026] = 1'b1; frame3.error[1026] = 1'b0;frame3.data[1027] = 8'hF8; frame3.valid[1027] = 1'b1; frame3.error[1027] = 1'b0;frame3.data[1028] = 8'hF9; frame3.valid[1028] = 1'b1; frame3.error[1028] = 1'b0;frame3.data[1029] = 8'hFA; frame3.valid[1029] = 1'b1; frame3.error[1029] = 1'b0;frame3.data[1030] = 8'hFB; frame3.valid[1030] = 1'b1; frame3.error[1030] = 1'b0;frame3.data[1031] = 8'hFC; frame3.valid[1031] = 1'b1; frame3.error[1031] = 1'b0;frame3.data[1032] = 8'hFD; frame3.valid[1032] = 1'b1; frame3.error[1032] = 1'b0;frame3.data[1033] = 8'hFE; frame3.valid[1033] = 1'b1; frame3.error[1033] = 1'b0;frame3.data[1034] = 8'h00; frame3.valid[1034] = 1'b1; frame3.error[1034] = 1'b0;frame3.data[1035] = 8'h01; frame3.valid[1035] = 1'b1; frame3.error[1035] = 1'b0;frame3.data[1036] = 8'h02; frame3.valid[1036] = 1'b1; frame3.error[1036] = 1'b0;frame3.data[1037] = 8'h03; frame3.valid[1037] = 1'b1; frame3.error[1037] = 1'b0;
        frame3.data[1038] = 8'h04; frame3.valid[1038] = 1'b1; frame3.error[1038] = 1'b0;frame3.data[1039] = 8'h05; frame3.valid[1039] = 1'b1; frame3.error[1039] = 1'b0;frame3.data[1040] = 8'h06; frame3.valid[1040] = 1'b1; frame3.error[1040] = 1'b0;frame3.data[1041] = 8'h07; frame3.valid[1041] = 1'b1; frame3.error[1041] = 1'b0;frame3.data[1042] = 8'h08; frame3.valid[1042] = 1'b1; frame3.error[1042] = 1'b0;frame3.data[1043] = 8'h09; frame3.valid[1043] = 1'b1; frame3.error[1043] = 1'b0;frame3.data[1044] = 8'h0A; frame3.valid[1044] = 1'b1; frame3.error[1044] = 1'b0;frame3.data[1045] = 8'h0B; frame3.valid[1045] = 1'b1; frame3.error[1045] = 1'b0;frame3.data[1046] = 8'h0C; frame3.valid[1046] = 1'b1; frame3.error[1046] = 1'b0;frame3.data[1047] = 8'h0D; frame3.valid[1047] = 1'b1; frame3.error[1047] = 1'b0;frame3.data[1048] = 8'h0E; frame3.valid[1048] = 1'b1; frame3.error[1048] = 1'b0;frame3.data[1049] = 8'h0F; frame3.valid[1049] = 1'b1; frame3.error[1049] = 1'b0;frame3.data[1050] = 8'h10; frame3.valid[1050] = 1'b1; frame3.error[1050] = 1'b0;frame3.data[1051] = 8'h11; frame3.valid[1051] = 1'b1; frame3.error[1051] = 1'b0;frame3.data[1052] = 8'h12; frame3.valid[1052] = 1'b1; frame3.error[1052] = 1'b0;frame3.data[1053] = 8'h13; frame3.valid[1053] = 1'b1; frame3.error[1053] = 1'b0;
        frame3.data[1054] = 8'h14; frame3.valid[1054] = 1'b1; frame3.error[1054] = 1'b0;frame3.data[1055] = 8'h15; frame3.valid[1055] = 1'b1; frame3.error[1055] = 1'b0;frame3.data[1056] = 8'h16; frame3.valid[1056] = 1'b1; frame3.error[1056] = 1'b0;frame3.data[1057] = 8'h17; frame3.valid[1057] = 1'b1; frame3.error[1057] = 1'b0;frame3.data[1058] = 8'h18; frame3.valid[1058] = 1'b1; frame3.error[1058] = 1'b0;frame3.data[1059] = 8'h19; frame3.valid[1059] = 1'b1; frame3.error[1059] = 1'b0;frame3.data[1060] = 8'h1A; frame3.valid[1060] = 1'b1; frame3.error[1060] = 1'b0;frame3.data[1061] = 8'h1B; frame3.valid[1061] = 1'b1; frame3.error[1061] = 1'b0;frame3.data[1062] = 8'h1C; frame3.valid[1062] = 1'b1; frame3.error[1062] = 1'b0;frame3.data[1063] = 8'h1D; frame3.valid[1063] = 1'b1; frame3.error[1063] = 1'b0;frame3.data[1064] = 8'h1E; frame3.valid[1064] = 1'b1; frame3.error[1064] = 1'b0;frame3.data[1065] = 8'h1F; frame3.valid[1065] = 1'b1; frame3.error[1065] = 1'b0;frame3.data[1066] = 8'h20; frame3.valid[1066] = 1'b1; frame3.error[1066] = 1'b0;frame3.data[1067] = 8'h21; frame3.valid[1067] = 1'b1; frame3.error[1067] = 1'b0;frame3.data[1068] = 8'h22; frame3.valid[1068] = 1'b1; frame3.error[1068] = 1'b0;frame3.data[1069] = 8'h23; frame3.valid[1069] = 1'b1; frame3.error[1069] = 1'b0;
        frame3.data[1070] = 8'h24; frame3.valid[1070] = 1'b1; frame3.error[1070] = 1'b0;frame3.data[1071] = 8'h25; frame3.valid[1071] = 1'b1; frame3.error[1071] = 1'b0;frame3.data[1072] = 8'h26; frame3.valid[1072] = 1'b1; frame3.error[1072] = 1'b0;frame3.data[1073] = 8'h27; frame3.valid[1073] = 1'b1; frame3.error[1073] = 1'b0;frame3.data[1074] = 8'h28; frame3.valid[1074] = 1'b1; frame3.error[1074] = 1'b0;frame3.data[1075] = 8'h29; frame3.valid[1075] = 1'b1; frame3.error[1075] = 1'b0;frame3.data[1076] = 8'h2A; frame3.valid[1076] = 1'b1; frame3.error[1076] = 1'b0;frame3.data[1077] = 8'h2B; frame3.valid[1077] = 1'b1; frame3.error[1077] = 1'b0;frame3.data[1078] = 8'h2C; frame3.valid[1078] = 1'b1; frame3.error[1078] = 1'b0;frame3.data[1079] = 8'h2D; frame3.valid[1079] = 1'b1; frame3.error[1079] = 1'b0;frame3.data[1080] = 8'h2E; frame3.valid[1080] = 1'b1; frame3.error[1080] = 1'b0;frame3.data[1081] = 8'h2F; frame3.valid[1081] = 1'b1; frame3.error[1081] = 1'b0;frame3.data[1082] = 8'h30; frame3.valid[1082] = 1'b1; frame3.error[1082] = 1'b0;frame3.data[1083] = 8'h31; frame3.valid[1083] = 1'b1; frame3.error[1083] = 1'b0;frame3.data[1084] = 8'h32; frame3.valid[1084] = 1'b1; frame3.error[1084] = 1'b0;frame3.data[1085] = 8'h33; frame3.valid[1085] = 1'b1; frame3.error[1085] = 1'b0;
        frame3.data[1086] = 8'h34; frame3.valid[1086] = 1'b1; frame3.error[1086] = 1'b0;frame3.data[1087] = 8'h35; frame3.valid[1087] = 1'b1; frame3.error[1087] = 1'b0;frame3.data[1088] = 8'h36; frame3.valid[1088] = 1'b1; frame3.error[1088] = 1'b0;frame3.data[1089] = 8'h37; frame3.valid[1089] = 1'b1; frame3.error[1089] = 1'b0;frame3.data[1090] = 8'h38; frame3.valid[1090] = 1'b1; frame3.error[1090] = 1'b0;frame3.data[1091] = 8'h39; frame3.valid[1091] = 1'b1; frame3.error[1091] = 1'b0;frame3.data[1092] = 8'h3A; frame3.valid[1092] = 1'b1; frame3.error[1092] = 1'b0;frame3.data[1093] = 8'h3B; frame3.valid[1093] = 1'b1; frame3.error[1093] = 1'b0;frame3.data[1094] = 8'h3C; frame3.valid[1094] = 1'b1; frame3.error[1094] = 1'b0;frame3.data[1095] = 8'h3D; frame3.valid[1095] = 1'b1; frame3.error[1095] = 1'b0;frame3.data[1096] = 8'h3E; frame3.valid[1096] = 1'b1; frame3.error[1096] = 1'b0;frame3.data[1097] = 8'h3F; frame3.valid[1097] = 1'b1; frame3.error[1097] = 1'b0;frame3.data[1098] = 8'h40; frame3.valid[1098] = 1'b1; frame3.error[1098] = 1'b0;frame3.data[1099] = 8'h41; frame3.valid[1099] = 1'b1; frame3.error[1099] = 1'b0;frame3.data[1100] = 8'h42; frame3.valid[1100] = 1'b1; frame3.error[1100] = 1'b0;frame3.data[1101] = 8'h43; frame3.valid[1101] = 1'b1; frame3.error[1101] = 1'b0;
        frame3.data[1102] = 8'h44; frame3.valid[1102] = 1'b1; frame3.error[1102] = 1'b0;frame3.data[1103] = 8'h45; frame3.valid[1103] = 1'b1; frame3.error[1103] = 1'b0;frame3.data[1104] = 8'h46; frame3.valid[1104] = 1'b1; frame3.error[1104] = 1'b0;frame3.data[1105] = 8'h47; frame3.valid[1105] = 1'b1; frame3.error[1105] = 1'b0;frame3.data[1106] = 8'h48; frame3.valid[1106] = 1'b1; frame3.error[1106] = 1'b0;frame3.data[1107] = 8'h49; frame3.valid[1107] = 1'b1; frame3.error[1107] = 1'b0;frame3.data[1108] = 8'h4A; frame3.valid[1108] = 1'b1; frame3.error[1108] = 1'b0;frame3.data[1109] = 8'h4B; frame3.valid[1109] = 1'b1; frame3.error[1109] = 1'b0;frame3.data[1110] = 8'h4C; frame3.valid[1110] = 1'b1; frame3.error[1110] = 1'b0;frame3.data[1111] = 8'h4D; frame3.valid[1111] = 1'b1; frame3.error[1111] = 1'b0;frame3.data[1112] = 8'h4E; frame3.valid[1112] = 1'b1; frame3.error[1112] = 1'b0;frame3.data[1113] = 8'h4F; frame3.valid[1113] = 1'b1; frame3.error[1113] = 1'b0;frame3.data[1114] = 8'h50; frame3.valid[1114] = 1'b1; frame3.error[1114] = 1'b0;frame3.data[1115] = 8'h51; frame3.valid[1115] = 1'b1; frame3.error[1115] = 1'b0;frame3.data[1116] = 8'h52; frame3.valid[1116] = 1'b1; frame3.error[1116] = 1'b0;frame3.data[1117] = 8'h53; frame3.valid[1117] = 1'b1; frame3.error[1117] = 1'b0;
        frame3.data[1118] = 8'h54; frame3.valid[1118] = 1'b1; frame3.error[1118] = 1'b0;frame3.data[1119] = 8'h55; frame3.valid[1119] = 1'b1; frame3.error[1119] = 1'b0;frame3.data[1120] = 8'h56; frame3.valid[1120] = 1'b1; frame3.error[1120] = 1'b0;frame3.data[1121] = 8'h57; frame3.valid[1121] = 1'b1; frame3.error[1121] = 1'b0;frame3.data[1122] = 8'h58; frame3.valid[1122] = 1'b1; frame3.error[1122] = 1'b0;frame3.data[1123] = 8'h59; frame3.valid[1123] = 1'b1; frame3.error[1123] = 1'b0;frame3.data[1124] = 8'h5A; frame3.valid[1124] = 1'b1; frame3.error[1124] = 1'b0;frame3.data[1125] = 8'h5B; frame3.valid[1125] = 1'b1; frame3.error[1125] = 1'b0;frame3.data[1126] = 8'h5C; frame3.valid[1126] = 1'b1; frame3.error[1126] = 1'b0;frame3.data[1127] = 8'h5D; frame3.valid[1127] = 1'b1; frame3.error[1127] = 1'b0;frame3.data[1128] = 8'h5E; frame3.valid[1128] = 1'b1; frame3.error[1128] = 1'b0;frame3.data[1129] = 8'h5F; frame3.valid[1129] = 1'b1; frame3.error[1129] = 1'b0;frame3.data[1130] = 8'h60; frame3.valid[1130] = 1'b1; frame3.error[1130] = 1'b0;frame3.data[1131] = 8'h61; frame3.valid[1131] = 1'b1; frame3.error[1131] = 1'b0;frame3.data[1132] = 8'h62; frame3.valid[1132] = 1'b1; frame3.error[1132] = 1'b0;frame3.data[1133] = 8'h63; frame3.valid[1133] = 1'b1; frame3.error[1133] = 1'b0;
        frame3.data[1134] = 8'h64; frame3.valid[1134] = 1'b1; frame3.error[1134] = 1'b0;frame3.data[1135] = 8'h65; frame3.valid[1135] = 1'b1; frame3.error[1135] = 1'b0;frame3.data[1136] = 8'h66; frame3.valid[1136] = 1'b1; frame3.error[1136] = 1'b0;frame3.data[1137] = 8'h67; frame3.valid[1137] = 1'b1; frame3.error[1137] = 1'b0;frame3.data[1138] = 8'h68; frame3.valid[1138] = 1'b1; frame3.error[1138] = 1'b0;frame3.data[1139] = 8'h69; frame3.valid[1139] = 1'b1; frame3.error[1139] = 1'b0;frame3.data[1140] = 8'h6A; frame3.valid[1140] = 1'b1; frame3.error[1140] = 1'b0;frame3.data[1141] = 8'h6B; frame3.valid[1141] = 1'b1; frame3.error[1141] = 1'b0;frame3.data[1142] = 8'h6C; frame3.valid[1142] = 1'b1; frame3.error[1142] = 1'b0;frame3.data[1143] = 8'h6D; frame3.valid[1143] = 1'b1; frame3.error[1143] = 1'b0;frame3.data[1144] = 8'h6E; frame3.valid[1144] = 1'b1; frame3.error[1144] = 1'b0;frame3.data[1145] = 8'h6F; frame3.valid[1145] = 1'b1; frame3.error[1145] = 1'b0;frame3.data[1146] = 8'h70; frame3.valid[1146] = 1'b1; frame3.error[1146] = 1'b0;frame3.data[1147] = 8'h71; frame3.valid[1147] = 1'b1; frame3.error[1147] = 1'b0;frame3.data[1148] = 8'h72; frame3.valid[1148] = 1'b1; frame3.error[1148] = 1'b0;frame3.data[1149] = 8'h73; frame3.valid[1149] = 1'b1; frame3.error[1149] = 1'b0;
        frame3.data[1150] = 8'h74; frame3.valid[1150] = 1'b1; frame3.error[1150] = 1'b0;frame3.data[1151] = 8'h75; frame3.valid[1151] = 1'b1; frame3.error[1151] = 1'b0;frame3.data[1152] = 8'h76; frame3.valid[1152] = 1'b1; frame3.error[1152] = 1'b0;frame3.data[1153] = 8'h77; frame3.valid[1153] = 1'b1; frame3.error[1153] = 1'b0;frame3.data[1154] = 8'h78; frame3.valid[1154] = 1'b1; frame3.error[1154] = 1'b0;frame3.data[1155] = 8'h79; frame3.valid[1155] = 1'b1; frame3.error[1155] = 1'b0;frame3.data[1156] = 8'h7A; frame3.valid[1156] = 1'b1; frame3.error[1156] = 1'b0;frame3.data[1157] = 8'h7B; frame3.valid[1157] = 1'b1; frame3.error[1157] = 1'b0;frame3.data[1158] = 8'h7C; frame3.valid[1158] = 1'b1; frame3.error[1158] = 1'b0;frame3.data[1159] = 8'h7D; frame3.valid[1159] = 1'b1; frame3.error[1159] = 1'b0;frame3.data[1160] = 8'h7E; frame3.valid[1160] = 1'b1; frame3.error[1160] = 1'b0;frame3.data[1161] = 8'h7F; frame3.valid[1161] = 1'b1; frame3.error[1161] = 1'b0;frame3.data[1162] = 8'h80; frame3.valid[1162] = 1'b1; frame3.error[1162] = 1'b0;frame3.data[1163] = 8'h81; frame3.valid[1163] = 1'b1; frame3.error[1163] = 1'b0;frame3.data[1164] = 8'h82; frame3.valid[1164] = 1'b1; frame3.error[1164] = 1'b0;frame3.data[1165] = 8'h83; frame3.valid[1165] = 1'b1; frame3.error[1165] = 1'b0;
        frame3.data[1166] = 8'h84; frame3.valid[1166] = 1'b1; frame3.error[1166] = 1'b0;frame3.data[1167] = 8'h85; frame3.valid[1167] = 1'b1; frame3.error[1167] = 1'b0;frame3.data[1168] = 8'h86; frame3.valid[1168] = 1'b1; frame3.error[1168] = 1'b0;frame3.data[1169] = 8'h87; frame3.valid[1169] = 1'b1; frame3.error[1169] = 1'b0;frame3.data[1170] = 8'h88; frame3.valid[1170] = 1'b1; frame3.error[1170] = 1'b0;frame3.data[1171] = 8'h89; frame3.valid[1171] = 1'b1; frame3.error[1171] = 1'b0;frame3.data[1172] = 8'h8A; frame3.valid[1172] = 1'b1; frame3.error[1172] = 1'b0;frame3.data[1173] = 8'h8B; frame3.valid[1173] = 1'b1; frame3.error[1173] = 1'b0;frame3.data[1174] = 8'h8C; frame3.valid[1174] = 1'b1; frame3.error[1174] = 1'b0;frame3.data[1175] = 8'h8D; frame3.valid[1175] = 1'b1; frame3.error[1175] = 1'b0;frame3.data[1176] = 8'h8E; frame3.valid[1176] = 1'b1; frame3.error[1176] = 1'b0;frame3.data[1177] = 8'h8F; frame3.valid[1177] = 1'b1; frame3.error[1177] = 1'b0;frame3.data[1178] = 8'h90; frame3.valid[1178] = 1'b1; frame3.error[1178] = 1'b0;frame3.data[1179] = 8'h91; frame3.valid[1179] = 1'b1; frame3.error[1179] = 1'b0;frame3.data[1180] = 8'h92; frame3.valid[1180] = 1'b1; frame3.error[1180] = 1'b0;frame3.data[1181] = 8'h93; frame3.valid[1181] = 1'b1; frame3.error[1181] = 1'b0;
        frame3.data[1182] = 8'h94; frame3.valid[1182] = 1'b1; frame3.error[1182] = 1'b0;frame3.data[1183] = 8'h95; frame3.valid[1183] = 1'b1; frame3.error[1183] = 1'b0;frame3.data[1184] = 8'h96; frame3.valid[1184] = 1'b1; frame3.error[1184] = 1'b0;frame3.data[1185] = 8'h97; frame3.valid[1185] = 1'b1; frame3.error[1185] = 1'b0;frame3.data[1186] = 8'h98; frame3.valid[1186] = 1'b1; frame3.error[1186] = 1'b0;frame3.data[1187] = 8'h99; frame3.valid[1187] = 1'b1; frame3.error[1187] = 1'b0;frame3.data[1188] = 8'h9A; frame3.valid[1188] = 1'b1; frame3.error[1188] = 1'b0;frame3.data[1189] = 8'h9B; frame3.valid[1189] = 1'b1; frame3.error[1189] = 1'b0;frame3.data[1190] = 8'h9C; frame3.valid[1190] = 1'b1; frame3.error[1190] = 1'b0;frame3.data[1191] = 8'h9D; frame3.valid[1191] = 1'b1; frame3.error[1191] = 1'b0;frame3.data[1192] = 8'h9E; frame3.valid[1192] = 1'b1; frame3.error[1192] = 1'b0;frame3.data[1193] = 8'h9F; frame3.valid[1193] = 1'b1; frame3.error[1193] = 1'b0;frame3.data[1194] = 8'hA0; frame3.valid[1194] = 1'b1; frame3.error[1194] = 1'b0;frame3.data[1195] = 8'hA1; frame3.valid[1195] = 1'b1; frame3.error[1195] = 1'b0;frame3.data[1196] = 8'hA2; frame3.valid[1196] = 1'b1; frame3.error[1196] = 1'b0;frame3.data[1197] = 8'hA3; frame3.valid[1197] = 1'b1; frame3.error[1197] = 1'b0;
        frame3.data[1198] = 8'hA4; frame3.valid[1198] = 1'b1; frame3.error[1198] = 1'b0;frame3.data[1199] = 8'hA5; frame3.valid[1199] = 1'b1; frame3.error[1199] = 1'b0;frame3.data[1200] = 8'hA6; frame3.valid[1200] = 1'b1; frame3.error[1200] = 1'b0;frame3.data[1201] = 8'hA7; frame3.valid[1201] = 1'b1; frame3.error[1201] = 1'b0;frame3.data[1202] = 8'hA8; frame3.valid[1202] = 1'b1; frame3.error[1202] = 1'b0;frame3.data[1203] = 8'hA9; frame3.valid[1203] = 1'b1; frame3.error[1203] = 1'b0;frame3.data[1204] = 8'hAA; frame3.valid[1204] = 1'b1; frame3.error[1204] = 1'b0;frame3.data[1205] = 8'hAB; frame3.valid[1205] = 1'b1; frame3.error[1205] = 1'b0;frame3.data[1206] = 8'hAC; frame3.valid[1206] = 1'b1; frame3.error[1206] = 1'b0;frame3.data[1207] = 8'hAD; frame3.valid[1207] = 1'b1; frame3.error[1207] = 1'b0;frame3.data[1208] = 8'hAE; frame3.valid[1208] = 1'b1; frame3.error[1208] = 1'b0;frame3.data[1209] = 8'hAF; frame3.valid[1209] = 1'b1; frame3.error[1209] = 1'b0;frame3.data[1210] = 8'hB0; frame3.valid[1210] = 1'b1; frame3.error[1210] = 1'b0;frame3.data[1211] = 8'hB1; frame3.valid[1211] = 1'b1; frame3.error[1211] = 1'b0;frame3.data[1212] = 8'hB2; frame3.valid[1212] = 1'b1; frame3.error[1212] = 1'b0;frame3.data[1213] = 8'hB3; frame3.valid[1213] = 1'b1; frame3.error[1213] = 1'b0;
        frame3.data[1214] = 8'hB4; frame3.valid[1214] = 1'b1; frame3.error[1214] = 1'b0;frame3.data[1215] = 8'hB5; frame3.valid[1215] = 1'b1; frame3.error[1215] = 1'b0;frame3.data[1216] = 8'hB6; frame3.valid[1216] = 1'b1; frame3.error[1216] = 1'b0;frame3.data[1217] = 8'hB7; frame3.valid[1217] = 1'b1; frame3.error[1217] = 1'b0;frame3.data[1218] = 8'hB8; frame3.valid[1218] = 1'b1; frame3.error[1218] = 1'b0;frame3.data[1219] = 8'hB9; frame3.valid[1219] = 1'b1; frame3.error[1219] = 1'b0;frame3.data[1220] = 8'hBA; frame3.valid[1220] = 1'b1; frame3.error[1220] = 1'b0;frame3.data[1221] = 8'hBB; frame3.valid[1221] = 1'b1; frame3.error[1221] = 1'b0;frame3.data[1222] = 8'hBC; frame3.valid[1222] = 1'b1; frame3.error[1222] = 1'b0;frame3.data[1223] = 8'hBD; frame3.valid[1223] = 1'b1; frame3.error[1223] = 1'b0;frame3.data[1224] = 8'hBE; frame3.valid[1224] = 1'b1; frame3.error[1224] = 1'b0;frame3.data[1225] = 8'hBF; frame3.valid[1225] = 1'b1; frame3.error[1225] = 1'b0;frame3.data[1226] = 8'hC0; frame3.valid[1226] = 1'b1; frame3.error[1226] = 1'b0;frame3.data[1227] = 8'hC1; frame3.valid[1227] = 1'b1; frame3.error[1227] = 1'b0;frame3.data[1228] = 8'hC2; frame3.valid[1228] = 1'b1; frame3.error[1228] = 1'b0;frame3.data[1229] = 8'hC3; frame3.valid[1229] = 1'b1; frame3.error[1229] = 1'b0;
        frame3.data[1230] = 8'hC4; frame3.valid[1230] = 1'b1; frame3.error[1230] = 1'b0;frame3.data[1231] = 8'hC5; frame3.valid[1231] = 1'b1; frame3.error[1231] = 1'b0;frame3.data[1232] = 8'hC6; frame3.valid[1232] = 1'b1; frame3.error[1232] = 1'b0;frame3.data[1233] = 8'hC7; frame3.valid[1233] = 1'b1; frame3.error[1233] = 1'b0;frame3.data[1234] = 8'hC8; frame3.valid[1234] = 1'b1; frame3.error[1234] = 1'b0;frame3.data[1235] = 8'hC9; frame3.valid[1235] = 1'b1; frame3.error[1235] = 1'b0;frame3.data[1236] = 8'hCA; frame3.valid[1236] = 1'b1; frame3.error[1236] = 1'b0;frame3.data[1237] = 8'hCB; frame3.valid[1237] = 1'b1; frame3.error[1237] = 1'b0;frame3.data[1238] = 8'hCC; frame3.valid[1238] = 1'b1; frame3.error[1238] = 1'b0;frame3.data[1239] = 8'hCD; frame3.valid[1239] = 1'b1; frame3.error[1239] = 1'b0;frame3.data[1240] = 8'hCE; frame3.valid[1240] = 1'b1; frame3.error[1240] = 1'b0;frame3.data[1241] = 8'hCF; frame3.valid[1241] = 1'b1; frame3.error[1241] = 1'b0;frame3.data[1242] = 8'hD0; frame3.valid[1242] = 1'b1; frame3.error[1242] = 1'b0;frame3.data[1243] = 8'hD1; frame3.valid[1243] = 1'b1; frame3.error[1243] = 1'b0;frame3.data[1244] = 8'hD2; frame3.valid[1244] = 1'b1; frame3.error[1244] = 1'b0;frame3.data[1245] = 8'hD3; frame3.valid[1245] = 1'b1; frame3.error[1245] = 1'b0;
        frame3.data[1246] = 8'hD4; frame3.valid[1246] = 1'b1; frame3.error[1246] = 1'b0;frame3.data[1247] = 8'hD5; frame3.valid[1247] = 1'b1; frame3.error[1247] = 1'b0;frame3.data[1248] = 8'hD6; frame3.valid[1248] = 1'b1; frame3.error[1248] = 1'b0;frame3.data[1249] = 8'hD7; frame3.valid[1249] = 1'b1; frame3.error[1249] = 1'b0;frame3.data[1250] = 8'hD8; frame3.valid[1250] = 1'b1; frame3.error[1250] = 1'b0;frame3.data[1251] = 8'hD9; frame3.valid[1251] = 1'b1; frame3.error[1251] = 1'b0;frame3.data[1252] = 8'hDA; frame3.valid[1252] = 1'b1; frame3.error[1252] = 1'b0;frame3.data[1253] = 8'hDB; frame3.valid[1253] = 1'b1; frame3.error[1253] = 1'b0;frame3.data[1254] = 8'hDC; frame3.valid[1254] = 1'b1; frame3.error[1254] = 1'b0;frame3.data[1255] = 8'hDD; frame3.valid[1255] = 1'b1; frame3.error[1255] = 1'b0;frame3.data[1256] = 8'hDE; frame3.valid[1256] = 1'b1; frame3.error[1256] = 1'b0;frame3.data[1257] = 8'hDF; frame3.valid[1257] = 1'b1; frame3.error[1257] = 1'b0;frame3.data[1258] = 8'hE0; frame3.valid[1258] = 1'b1; frame3.error[1258] = 1'b0;frame3.data[1259] = 8'hE1; frame3.valid[1259] = 1'b1; frame3.error[1259] = 1'b0;frame3.data[1260] = 8'hE2; frame3.valid[1260] = 1'b1; frame3.error[1260] = 1'b0;frame3.data[1261] = 8'hE3; frame3.valid[1261] = 1'b1; frame3.error[1261] = 1'b0;
        frame3.data[1262] = 8'hE4; frame3.valid[1262] = 1'b1; frame3.error[1262] = 1'b0;frame3.data[1263] = 8'hE5; frame3.valid[1263] = 1'b1; frame3.error[1263] = 1'b0;frame3.data[1264] = 8'hE6; frame3.valid[1264] = 1'b1; frame3.error[1264] = 1'b0;frame3.data[1265] = 8'hE7; frame3.valid[1265] = 1'b1; frame3.error[1265] = 1'b0;frame3.data[1266] = 8'hE8; frame3.valid[1266] = 1'b1; frame3.error[1266] = 1'b0;frame3.data[1267] = 8'hE9; frame3.valid[1267] = 1'b1; frame3.error[1267] = 1'b0;frame3.data[1268] = 8'hEA; frame3.valid[1268] = 1'b1; frame3.error[1268] = 1'b0;frame3.data[1269] = 8'hEB; frame3.valid[1269] = 1'b1; frame3.error[1269] = 1'b0;frame3.data[1270] = 8'hEC; frame3.valid[1270] = 1'b1; frame3.error[1270] = 1'b0;frame3.data[1271] = 8'hED; frame3.valid[1271] = 1'b1; frame3.error[1271] = 1'b0;frame3.data[1272] = 8'hEE; frame3.valid[1272] = 1'b1; frame3.error[1272] = 1'b0;frame3.data[1273] = 8'hEF; frame3.valid[1273] = 1'b1; frame3.error[1273] = 1'b0;frame3.data[1274] = 8'hF0; frame3.valid[1274] = 1'b1; frame3.error[1274] = 1'b0;frame3.data[1275] = 8'hF1; frame3.valid[1275] = 1'b1; frame3.error[1275] = 1'b0;frame3.data[1276] = 8'hF2; frame3.valid[1276] = 1'b1; frame3.error[1276] = 1'b0;frame3.data[1277] = 8'hF3; frame3.valid[1277] = 1'b1; frame3.error[1277] = 1'b0;
        frame3.data[1278] = 8'hF4; frame3.valid[1278] = 1'b1; frame3.error[1278] = 1'b0;frame3.data[1279] = 8'hF5; frame3.valid[1279] = 1'b1; frame3.error[1279] = 1'b0;frame3.data[1280] = 8'hF6; frame3.valid[1280] = 1'b1; frame3.error[1280] = 1'b0;frame3.data[1281] = 8'hF7; frame3.valid[1281] = 1'b1; frame3.error[1281] = 1'b0;frame3.data[1282] = 8'hF8; frame3.valid[1282] = 1'b1; frame3.error[1282] = 1'b0;frame3.data[1283] = 8'hF9; frame3.valid[1283] = 1'b1; frame3.error[1283] = 1'b0;frame3.data[1284] = 8'hFA; frame3.valid[1284] = 1'b1; frame3.error[1284] = 1'b0;frame3.data[1285] = 8'hFB; frame3.valid[1285] = 1'b1; frame3.error[1285] = 1'b0;frame3.data[1286] = 8'hFC; frame3.valid[1286] = 1'b1; frame3.error[1286] = 1'b0;frame3.data[1287] = 8'hFD; frame3.valid[1287] = 1'b1; frame3.error[1287] = 1'b0;frame3.data[1288] = 8'hFE; frame3.valid[1288] = 1'b1; frame3.error[1288] = 1'b0;frame3.data[1289] = 8'h00; frame3.valid[1289] = 1'b1; frame3.error[1289] = 1'b0;frame3.data[1290] = 8'h01; frame3.valid[1290] = 1'b1; frame3.error[1290] = 1'b0;frame3.data[1291] = 8'h02; frame3.valid[1291] = 1'b1; frame3.error[1291] = 1'b0;frame3.data[1292] = 8'h03; frame3.valid[1292] = 1'b1; frame3.error[1292] = 1'b0;frame3.data[1293] = 8'h04; frame3.valid[1293] = 1'b1; frame3.error[1293] = 1'b0;
        frame3.data[1294] = 8'h05; frame3.valid[1294] = 1'b1; frame3.error[1294] = 1'b0;frame3.data[1295] = 8'h06; frame3.valid[1295] = 1'b1; frame3.error[1295] = 1'b0;frame3.data[1296] = 8'h07; frame3.valid[1296] = 1'b1; frame3.error[1296] = 1'b0;frame3.data[1297] = 8'h08; frame3.valid[1297] = 1'b1; frame3.error[1297] = 1'b0;frame3.data[1298] = 8'h09; frame3.valid[1298] = 1'b1; frame3.error[1298] = 1'b0;frame3.data[1299] = 8'h0A; frame3.valid[1299] = 1'b1; frame3.error[1299] = 1'b0;frame3.data[1300] = 8'h0B; frame3.valid[1300] = 1'b1; frame3.error[1300] = 1'b0;frame3.data[1301] = 8'h0C; frame3.valid[1301] = 1'b1; frame3.error[1301] = 1'b0;frame3.data[1302] = 8'h0D; frame3.valid[1302] = 1'b1; frame3.error[1302] = 1'b0;frame3.data[1303] = 8'h0E; frame3.valid[1303] = 1'b1; frame3.error[1303] = 1'b0;frame3.data[1304] = 8'h0F; frame3.valid[1304] = 1'b1; frame3.error[1304] = 1'b0;frame3.data[1305] = 8'h10; frame3.valid[1305] = 1'b1; frame3.error[1305] = 1'b0;frame3.data[1306] = 8'h11; frame3.valid[1306] = 1'b1; frame3.error[1306] = 1'b0;frame3.data[1307] = 8'h12; frame3.valid[1307] = 1'b1; frame3.error[1307] = 1'b0;frame3.data[1308] = 8'h13; frame3.valid[1308] = 1'b1; frame3.error[1308] = 1'b0;frame3.data[1309] = 8'h14; frame3.valid[1309] = 1'b1; frame3.error[1309] = 1'b0;
        frame3.data[1310] = 8'h15; frame3.valid[1310] = 1'b1; frame3.error[1310] = 1'b0;frame3.data[1311] = 8'h16; frame3.valid[1311] = 1'b1; frame3.error[1311] = 1'b0;frame3.data[1312] = 8'h17; frame3.valid[1312] = 1'b1; frame3.error[1312] = 1'b0;frame3.data[1313] = 8'h18; frame3.valid[1313] = 1'b1; frame3.error[1313] = 1'b0;frame3.data[1314] = 8'h19; frame3.valid[1314] = 1'b1; frame3.error[1314] = 1'b0;frame3.data[1315] = 8'h1A; frame3.valid[1315] = 1'b1; frame3.error[1315] = 1'b0;frame3.data[1316] = 8'h1B; frame3.valid[1316] = 1'b1; frame3.error[1316] = 1'b0;frame3.data[1317] = 8'h1C; frame3.valid[1317] = 1'b1; frame3.error[1317] = 1'b0;frame3.data[1318] = 8'h1D; frame3.valid[1318] = 1'b1; frame3.error[1318] = 1'b0;frame3.data[1319] = 8'h1E; frame3.valid[1319] = 1'b1; frame3.error[1319] = 1'b0;frame3.data[1320] = 8'h1F; frame3.valid[1320] = 1'b1; frame3.error[1320] = 1'b0;frame3.data[1321] = 8'h20; frame3.valid[1321] = 1'b1; frame3.error[1321] = 1'b0;frame3.data[1322] = 8'h21; frame3.valid[1322] = 1'b1; frame3.error[1322] = 1'b0;frame3.data[1323] = 8'h22; frame3.valid[1323] = 1'b1; frame3.error[1323] = 1'b0;frame3.data[1324] = 8'h23; frame3.valid[1324] = 1'b1; frame3.error[1324] = 1'b0;frame3.data[1325] = 8'h24; frame3.valid[1325] = 1'b1; frame3.error[1325] = 1'b0;
        frame3.data[1326] = 8'h25; frame3.valid[1326] = 1'b1; frame3.error[1326] = 1'b0;frame3.data[1327] = 8'h26; frame3.valid[1327] = 1'b1; frame3.error[1327] = 1'b0;frame3.data[1328] = 8'h27; frame3.valid[1328] = 1'b1; frame3.error[1328] = 1'b0;frame3.data[1329] = 8'h28; frame3.valid[1329] = 1'b1; frame3.error[1329] = 1'b0;frame3.data[1330] = 8'h29; frame3.valid[1330] = 1'b1; frame3.error[1330] = 1'b0;frame3.data[1331] = 8'h2A; frame3.valid[1331] = 1'b1; frame3.error[1331] = 1'b0;frame3.data[1332] = 8'h2B; frame3.valid[1332] = 1'b1; frame3.error[1332] = 1'b0;frame3.data[1333] = 8'h2C; frame3.valid[1333] = 1'b1; frame3.error[1333] = 1'b0;frame3.data[1334] = 8'h2D; frame3.valid[1334] = 1'b1; frame3.error[1334] = 1'b0;frame3.data[1335] = 8'h2E; frame3.valid[1335] = 1'b1; frame3.error[1335] = 1'b0;frame3.data[1336] = 8'h2F; frame3.valid[1336] = 1'b1; frame3.error[1336] = 1'b0;frame3.data[1337] = 8'h30; frame3.valid[1337] = 1'b1; frame3.error[1337] = 1'b0;frame3.data[1338] = 8'h31; frame3.valid[1338] = 1'b1; frame3.error[1338] = 1'b0;frame3.data[1339] = 8'h32; frame3.valid[1339] = 1'b1; frame3.error[1339] = 1'b0;frame3.data[1340] = 8'h33; frame3.valid[1340] = 1'b1; frame3.error[1340] = 1'b0;frame3.data[1341] = 8'h34; frame3.valid[1341] = 1'b1; frame3.error[1341] = 1'b0;
        frame3.data[1342] = 8'h35; frame3.valid[1342] = 1'b1; frame3.error[1342] = 1'b0;frame3.data[1343] = 8'h36; frame3.valid[1343] = 1'b1; frame3.error[1343] = 1'b0;frame3.data[1344] = 8'h37; frame3.valid[1344] = 1'b1; frame3.error[1344] = 1'b0;frame3.data[1345] = 8'h38; frame3.valid[1345] = 1'b1; frame3.error[1345] = 1'b0;frame3.data[1346] = 8'h39; frame3.valid[1346] = 1'b1; frame3.error[1346] = 1'b0;frame3.data[1347] = 8'h3A; frame3.valid[1347] = 1'b1; frame3.error[1347] = 1'b0;frame3.data[1348] = 8'h3B; frame3.valid[1348] = 1'b1; frame3.error[1348] = 1'b0;frame3.data[1349] = 8'h3C; frame3.valid[1349] = 1'b1; frame3.error[1349] = 1'b0;frame3.data[1350] = 8'h3D; frame3.valid[1350] = 1'b1; frame3.error[1350] = 1'b0;frame3.data[1351] = 8'h3E; frame3.valid[1351] = 1'b1; frame3.error[1351] = 1'b0;frame3.data[1352] = 8'h3F; frame3.valid[1352] = 1'b1; frame3.error[1352] = 1'b0;frame3.data[1353] = 8'h40; frame3.valid[1353] = 1'b1; frame3.error[1353] = 1'b0;frame3.data[1354] = 8'h41; frame3.valid[1354] = 1'b1; frame3.error[1354] = 1'b0;frame3.data[1355] = 8'h42; frame3.valid[1355] = 1'b1; frame3.error[1355] = 1'b0;frame3.data[1356] = 8'h43; frame3.valid[1356] = 1'b1; frame3.error[1356] = 1'b0;frame3.data[1357] = 8'h44; frame3.valid[1357] = 1'b1; frame3.error[1357] = 1'b0;
        frame3.data[1358] = 8'h45; frame3.valid[1358] = 1'b1; frame3.error[1358] = 1'b0;frame3.data[1359] = 8'h46; frame3.valid[1359] = 1'b1; frame3.error[1359] = 1'b0;frame3.data[1360] = 8'h47; frame3.valid[1360] = 1'b1; frame3.error[1360] = 1'b0;frame3.data[1361] = 8'h48; frame3.valid[1361] = 1'b1; frame3.error[1361] = 1'b0;frame3.data[1362] = 8'h49; frame3.valid[1362] = 1'b1; frame3.error[1362] = 1'b0;frame3.data[1363] = 8'h4A; frame3.valid[1363] = 1'b1; frame3.error[1363] = 1'b0;frame3.data[1364] = 8'h4B; frame3.valid[1364] = 1'b1; frame3.error[1364] = 1'b0;frame3.data[1365] = 8'h4C; frame3.valid[1365] = 1'b1; frame3.error[1365] = 1'b0;frame3.data[1366] = 8'h4D; frame3.valid[1366] = 1'b1; frame3.error[1366] = 1'b0;frame3.data[1367] = 8'h4E; frame3.valid[1367] = 1'b1; frame3.error[1367] = 1'b0;frame3.data[1368] = 8'h4F; frame3.valid[1368] = 1'b1; frame3.error[1368] = 1'b0;frame3.data[1369] = 8'h50; frame3.valid[1369] = 1'b1; frame3.error[1369] = 1'b0;frame3.data[1370] = 8'h51; frame3.valid[1370] = 1'b1; frame3.error[1370] = 1'b0;frame3.data[1371] = 8'h52; frame3.valid[1371] = 1'b1; frame3.error[1371] = 1'b0;frame3.data[1372] = 8'h53; frame3.valid[1372] = 1'b1; frame3.error[1372] = 1'b0;frame3.data[1373] = 8'h54; frame3.valid[1373] = 1'b1; frame3.error[1373] = 1'b0;
        frame3.data[1374] = 8'h55; frame3.valid[1374] = 1'b1; frame3.error[1374] = 1'b0;frame3.data[1375] = 8'h56; frame3.valid[1375] = 1'b1; frame3.error[1375] = 1'b0;frame3.data[1376] = 8'h57; frame3.valid[1376] = 1'b1; frame3.error[1376] = 1'b0;frame3.data[1377] = 8'h58; frame3.valid[1377] = 1'b1; frame3.error[1377] = 1'b0;frame3.data[1378] = 8'h59; frame3.valid[1378] = 1'b1; frame3.error[1378] = 1'b0;frame3.data[1379] = 8'h5A; frame3.valid[1379] = 1'b1; frame3.error[1379] = 1'b0;frame3.data[1380] = 8'h5B; frame3.valid[1380] = 1'b1; frame3.error[1380] = 1'b0;frame3.data[1381] = 8'h5C; frame3.valid[1381] = 1'b1; frame3.error[1381] = 1'b0;frame3.data[1382] = 8'h5D; frame3.valid[1382] = 1'b1; frame3.error[1382] = 1'b0;frame3.data[1383] = 8'h5E; frame3.valid[1383] = 1'b1; frame3.error[1383] = 1'b0;frame3.data[1384] = 8'h5F; frame3.valid[1384] = 1'b1; frame3.error[1384] = 1'b0;frame3.data[1385] = 8'h60; frame3.valid[1385] = 1'b1; frame3.error[1385] = 1'b0;frame3.data[1386] = 8'h61; frame3.valid[1386] = 1'b1; frame3.error[1386] = 1'b0;frame3.data[1387] = 8'h62; frame3.valid[1387] = 1'b1; frame3.error[1387] = 1'b0;frame3.data[1388] = 8'h63; frame3.valid[1388] = 1'b1; frame3.error[1388] = 1'b0;frame3.data[1389] = 8'h64; frame3.valid[1389] = 1'b1; frame3.error[1389] = 1'b0;
        frame3.data[1390] = 8'h65; frame3.valid[1390] = 1'b1; frame3.error[1390] = 1'b0;frame3.data[1391] = 8'h66; frame3.valid[1391] = 1'b1; frame3.error[1391] = 1'b0;frame3.data[1392] = 8'h67; frame3.valid[1392] = 1'b1; frame3.error[1392] = 1'b0;frame3.data[1393] = 8'h68; frame3.valid[1393] = 1'b1; frame3.error[1393] = 1'b0;frame3.data[1394] = 8'h69; frame3.valid[1394] = 1'b1; frame3.error[1394] = 1'b0;frame3.data[1395] = 8'h6A; frame3.valid[1395] = 1'b1; frame3.error[1395] = 1'b0;frame3.data[1396] = 8'h6B; frame3.valid[1396] = 1'b1; frame3.error[1396] = 1'b0;frame3.data[1397] = 8'h6C; frame3.valid[1397] = 1'b1; frame3.error[1397] = 1'b0;frame3.data[1398] = 8'h6D; frame3.valid[1398] = 1'b1; frame3.error[1398] = 1'b0;frame3.data[1399] = 8'h6E; frame3.valid[1399] = 1'b1; frame3.error[1399] = 1'b0;frame3.data[1400] = 8'h6F; frame3.valid[1400] = 1'b1; frame3.error[1400] = 1'b0;frame3.data[1401] = 8'h70; frame3.valid[1401] = 1'b1; frame3.error[1401] = 1'b0;frame3.data[1402] = 8'h71; frame3.valid[1402] = 1'b1; frame3.error[1402] = 1'b0;frame3.data[1403] = 8'h72; frame3.valid[1403] = 1'b1; frame3.error[1403] = 1'b0;frame3.data[1404] = 8'h73; frame3.valid[1404] = 1'b1; frame3.error[1404] = 1'b0;frame3.data[1405] = 8'h74; frame3.valid[1405] = 1'b1; frame3.error[1405] = 1'b0;
        frame3.data[1406] = 8'h75; frame3.valid[1406] = 1'b1; frame3.error[1406] = 1'b0;frame3.data[1407] = 8'h76; frame3.valid[1407] = 1'b1; frame3.error[1407] = 1'b0;frame3.data[1408] = 8'h77; frame3.valid[1408] = 1'b1; frame3.error[1408] = 1'b0;frame3.data[1409] = 8'h78; frame3.valid[1409] = 1'b1; frame3.error[1409] = 1'b0;frame3.data[1410] = 8'h79; frame3.valid[1410] = 1'b1; frame3.error[1410] = 1'b0;frame3.data[1411] = 8'h7A; frame3.valid[1411] = 1'b1; frame3.error[1411] = 1'b0;frame3.data[1412] = 8'h7B; frame3.valid[1412] = 1'b1; frame3.error[1412] = 1'b0;frame3.data[1413] = 8'h7C; frame3.valid[1413] = 1'b1; frame3.error[1413] = 1'b0;frame3.data[1414] = 8'h7D; frame3.valid[1414] = 1'b1; frame3.error[1414] = 1'b0;frame3.data[1415] = 8'h7E; frame3.valid[1415] = 1'b1; frame3.error[1415] = 1'b0;frame3.data[1416] = 8'h7F; frame3.valid[1416] = 1'b1; frame3.error[1416] = 1'b0;frame3.data[1417] = 8'h80; frame3.valid[1417] = 1'b1; frame3.error[1417] = 1'b0;frame3.data[1418] = 8'h81; frame3.valid[1418] = 1'b1; frame3.error[1418] = 1'b0;frame3.data[1419] = 8'h82; frame3.valid[1419] = 1'b1; frame3.error[1419] = 1'b0;frame3.data[1420] = 8'h83; frame3.valid[1420] = 1'b1; frame3.error[1420] = 1'b0;frame3.data[1421] = 8'h84; frame3.valid[1421] = 1'b1; frame3.error[1421] = 1'b0;
        frame3.data[1422] = 8'h85; frame3.valid[1422] = 1'b1; frame3.error[1422] = 1'b0;frame3.data[1423] = 8'h86; frame3.valid[1423] = 1'b1; frame3.error[1423] = 1'b0;frame3.data[1424] = 8'h87; frame3.valid[1424] = 1'b1; frame3.error[1424] = 1'b0;frame3.data[1425] = 8'h88; frame3.valid[1425] = 1'b1; frame3.error[1425] = 1'b0;frame3.data[1426] = 8'h89; frame3.valid[1426] = 1'b1; frame3.error[1426] = 1'b0;frame3.data[1427] = 8'h8A; frame3.valid[1427] = 1'b1; frame3.error[1427] = 1'b0;frame3.data[1428] = 8'h8B; frame3.valid[1428] = 1'b1; frame3.error[1428] = 1'b0;frame3.data[1429] = 8'h8C; frame3.valid[1429] = 1'b1; frame3.error[1429] = 1'b0;frame3.data[1430] = 8'h8D; frame3.valid[1430] = 1'b1; frame3.error[1430] = 1'b0;frame3.data[1431] = 8'h8E; frame3.valid[1431] = 1'b1; frame3.error[1431] = 1'b0;frame3.data[1432] = 8'h8F; frame3.valid[1432] = 1'b1; frame3.error[1432] = 1'b0;frame3.data[1433] = 8'h90; frame3.valid[1433] = 1'b1; frame3.error[1433] = 1'b0;frame3.data[1434] = 8'h91; frame3.valid[1434] = 1'b1; frame3.error[1434] = 1'b0;frame3.data[1435] = 8'h92; frame3.valid[1435] = 1'b1; frame3.error[1435] = 1'b0;frame3.data[1436] = 8'h93; frame3.valid[1436] = 1'b1; frame3.error[1436] = 1'b0;frame3.data[1437] = 8'h94; frame3.valid[1437] = 1'b1; frame3.error[1437] = 1'b0;
        frame3.data[1438] = 8'h95; frame3.valid[1438] = 1'b1; frame3.error[1438] = 1'b0;frame3.data[1439] = 8'h96; frame3.valid[1439] = 1'b1; frame3.error[1439] = 1'b0;frame3.data[1440] = 8'h97; frame3.valid[1440] = 1'b1; frame3.error[1440] = 1'b0;frame3.data[1441] = 8'h98; frame3.valid[1441] = 1'b1; frame3.error[1441] = 1'b0;frame3.data[1442] = 8'h99; frame3.valid[1442] = 1'b1; frame3.error[1442] = 1'b0;frame3.data[1443] = 8'h9A; frame3.valid[1443] = 1'b1; frame3.error[1443] = 1'b0;frame3.data[1444] = 8'h9B; frame3.valid[1444] = 1'b1; frame3.error[1444] = 1'b0;frame3.data[1445] = 8'h9C; frame3.valid[1445] = 1'b1; frame3.error[1445] = 1'b0;frame3.data[1446] = 8'h9D; frame3.valid[1446] = 1'b1; frame3.error[1446] = 1'b0;frame3.data[1447] = 8'h9E; frame3.valid[1447] = 1'b1; frame3.error[1447] = 1'b0;frame3.data[1448] = 8'h9F; frame3.valid[1448] = 1'b1; frame3.error[1448] = 1'b0;frame3.data[1449] = 8'hA0; frame3.valid[1449] = 1'b1; frame3.error[1449] = 1'b0;frame3.data[1450] = 8'hA1; frame3.valid[1450] = 1'b1; frame3.error[1450] = 1'b0;frame3.data[1451] = 8'hA2; frame3.valid[1451] = 1'b1; frame3.error[1451] = 1'b0;frame3.data[1452] = 8'hA3; frame3.valid[1452] = 1'b1; frame3.error[1452] = 1'b0;frame3.data[1453] = 8'hA4; frame3.valid[1453] = 1'b1; frame3.error[1453] = 1'b0;
        frame3.data[1454] = 8'hA5; frame3.valid[1454] = 1'b1; frame3.error[1454] = 1'b0;frame3.data[1455] = 8'hA6; frame3.valid[1455] = 1'b1; frame3.error[1455] = 1'b0;frame3.data[1456] = 8'hA7; frame3.valid[1456] = 1'b1; frame3.error[1456] = 1'b0;frame3.data[1457] = 8'hA8; frame3.valid[1457] = 1'b1; frame3.error[1457] = 1'b0;frame3.data[1458] = 8'hA9; frame3.valid[1458] = 1'b1; frame3.error[1458] = 1'b0;frame3.data[1459] = 8'hAA; frame3.valid[1459] = 1'b1; frame3.error[1459] = 1'b0;frame3.data[1460] = 8'hAB; frame3.valid[1460] = 1'b1; frame3.error[1460] = 1'b0;frame3.data[1461] = 8'hAC; frame3.valid[1461] = 1'b1; frame3.error[1461] = 1'b0;frame3.data[1462] = 8'hAD; frame3.valid[1462] = 1'b1; frame3.error[1462] = 1'b0;frame3.data[1463] = 8'hAE; frame3.valid[1463] = 1'b1; frame3.error[1463] = 1'b0;frame3.data[1464] = 8'hAF; frame3.valid[1464] = 1'b1; frame3.error[1464] = 1'b0;frame3.data[1465] = 8'hB0; frame3.valid[1465] = 1'b1; frame3.error[1465] = 1'b0;frame3.data[1466] = 8'hB1; frame3.valid[1466] = 1'b1; frame3.error[1466] = 1'b0;frame3.data[1467] = 8'hB2; frame3.valid[1467] = 1'b1; frame3.error[1467] = 1'b0;frame3.data[1468] = 8'hB3; frame3.valid[1468] = 1'b1; frame3.error[1468] = 1'b0;frame3.data[1469] = 8'hB4; frame3.valid[1469] = 1'b1; frame3.error[1469] = 1'b0;
        frame3.data[1470] = 8'hB5; frame3.valid[1470] = 1'b1; frame3.error[1470] = 1'b0;frame3.data[1471] = 8'hB6; frame3.valid[1471] = 1'b1; frame3.error[1471] = 1'b0;frame3.data[1472] = 8'hB7; frame3.valid[1472] = 1'b1; frame3.error[1472] = 1'b0;frame3.data[1473] = 8'hB8; frame3.valid[1473] = 1'b1; frame3.error[1473] = 1'b0;frame3.data[1474] = 8'hB9; frame3.valid[1474] = 1'b1; frame3.error[1474] = 1'b0;frame3.data[1475] = 8'hBA; frame3.valid[1475] = 1'b1; frame3.error[1475] = 1'b0;frame3.data[1476] = 8'hBB; frame3.valid[1476] = 1'b1; frame3.error[1476] = 1'b0;frame3.data[1477] = 8'hBC; frame3.valid[1477] = 1'b1; frame3.error[1477] = 1'b0;frame3.data[1478] = 8'hBD; frame3.valid[1478] = 1'b1; frame3.error[1478] = 1'b0;frame3.data[1479] = 8'hBE; frame3.valid[1479] = 1'b1; frame3.error[1479] = 1'b0;frame3.data[1480] = 8'hBF; frame3.valid[1480] = 1'b1; frame3.error[1480] = 1'b0;frame3.data[1481] = 8'hC0; frame3.valid[1481] = 1'b1; frame3.error[1481] = 1'b0;frame3.data[1482] = 8'hC1; frame3.valid[1482] = 1'b1; frame3.error[1482] = 1'b0;frame3.data[1483] = 8'hC2; frame3.valid[1483] = 1'b1; frame3.error[1483] = 1'b0;frame3.data[1484] = 8'hC3; frame3.valid[1484] = 1'b1; frame3.error[1484] = 1'b0;frame3.data[1485] = 8'hC4; frame3.valid[1485] = 1'b1; frame3.error[1485] = 1'b0;
        frame3.data[1486] = 8'hC5; frame3.valid[1486] = 1'b1; frame3.error[1486] = 1'b0;frame3.data[1487] = 8'hC6; frame3.valid[1487] = 1'b1; frame3.error[1487] = 1'b0;frame3.data[1488] = 8'hC7; frame3.valid[1488] = 1'b1; frame3.error[1488] = 1'b0;frame3.data[1489] = 8'hC8; frame3.valid[1489] = 1'b1; frame3.error[1489] = 1'b0;frame3.data[1490] = 8'hC9; frame3.valid[1490] = 1'b1; frame3.error[1490] = 1'b0;frame3.data[1491] = 8'hCA; frame3.valid[1491] = 1'b1; frame3.error[1491] = 1'b0;frame3.data[1492] = 8'hCB; frame3.valid[1492] = 1'b1; frame3.error[1492] = 1'b0;frame3.data[1493] = 8'hCC; frame3.valid[1493] = 1'b1; frame3.error[1493] = 1'b0;frame3.data[1494] = 8'hCD; frame3.valid[1494] = 1'b1; frame3.error[1494] = 1'b0;frame3.data[1495] = 8'hCE; frame3.valid[1495] = 1'b1; frame3.error[1495] = 1'b0;frame3.data[1496] = 8'hCF; frame3.valid[1496] = 1'b1; frame3.error[1496] = 1'b0;frame3.data[1497] = 8'hD0; frame3.valid[1497] = 1'b1; frame3.error[1497] = 1'b0;frame3.data[1498] = 8'hD1; frame3.valid[1498] = 1'b1; frame3.error[1498] = 1'b0;frame3.data[1499] = 8'hD2; frame3.valid[1499] = 1'b1; frame3.error[1499] = 1'b0;frame3.data[1500] = 8'hD3; frame3.valid[1500] = 1'b1; frame3.error[1500] = 1'b0;frame3.data[1501] = 8'hD4; frame3.valid[1501] = 1'b1; frame3.error[1501] = 1'b0;
        frame3.data[1502] = 8'hD5; frame3.valid[1502] = 1'b1; frame3.error[1502] = 1'b0;frame3.data[1503] = 8'hD6; frame3.valid[1503] = 1'b1; frame3.error[1503] = 1'b0;frame3.data[1504] = 8'hD7; frame3.valid[1504] = 1'b1; frame3.error[1504] = 1'b0;frame3.data[1505] = 8'hD8; frame3.valid[1505] = 1'b1; frame3.error[1505] = 1'b0;frame3.data[1506] = 8'hD9; frame3.valid[1506] = 1'b1; frame3.error[1506] = 1'b0;frame3.data[1507] = 8'hDA; frame3.valid[1507] = 1'b1; frame3.error[1507] = 1'b0;frame3.data[1508] = 8'hDB; frame3.valid[1508] = 1'b1; frame3.error[1508] = 1'b0;frame3.data[1509] = 8'hDC; frame3.valid[1509] = 1'b1; frame3.error[1509] = 1'b0;frame3.data[1510] = 8'hDD; frame3.valid[1510] = 1'b1; frame3.error[1510] = 1'b0;frame3.data[1511] = 8'hDE; frame3.valid[1511] = 1'b1; frame3.error[1511] = 1'b0;frame3.data[1512] = 8'hDF; frame3.valid[1512] = 1'b1; frame3.error[1512] = 1'b0;frame3.data[1513] = 8'hE0; frame3.valid[1513] = 1'b1; frame3.error[1513] = 1'b0;


        frame3.data[1514] = 8'h00;  frame3.valid[1514] = 1'b0;  frame3.error[1514] = 1'b0;
        frame3.data[1515] = 8'h00;  frame3.valid[1515] = 1'b0;  frame3.error[1515] = 1'b0;

        // No error in this frame
        frame3.bad_frame  = 1'b0;

        payload_length = FRAME_LENGTH - 14;
        // {frame0.data[12], frame0.data[13]} = payload_length;
        // {frame1.data[12], frame1.data[13]} = payload_length;
        {frame2.data[12], frame2.data[13]} = payload_length;
        {frame3.data[12], frame3.data[13]} = payload_length;
        frame0.valid[FRAME_LENGTH] = 1'b0;
        frame1.valid[FRAME_LENGTH] = 1'b0;
        frame2.valid[FRAME_LENGTH] = 1'b0;
        frame3.valid[FRAME_LENGTH] = 1'b0;
    end

    //--------------------------------------------------------------------
    // CRC engine
    //--------------------------------------------------------------------
    task calc_crc;
        input  [7:0]  data;
        inout  [31:0] fcs;

        reg [31:0] crc;
        reg        crc_feedback;
        integer    I;
    begin

        crc = ~ fcs;

        for (I = 0; I < 8; I = I + 1)
        begin
            crc_feedback = crc[0] ^ data[I];

            crc[0]       = crc[1];
            crc[1]       = crc[2];
            crc[2]       = crc[3];
            crc[3]       = crc[4];
            crc[4]       = crc[5];
            crc[5]       = crc[6]  ^ crc_feedback;
            crc[6]       = crc[7];
            crc[7]       = crc[8];
            crc[8]       = crc[9]  ^ crc_feedback;
            crc[9]       = crc[10] ^ crc_feedback;
            crc[10]      = crc[11];
            crc[11]      = crc[12];
            crc[12]      = crc[13];
            crc[13]      = crc[14];
            crc[14]      = crc[15];
            crc[15]      = crc[16] ^ crc_feedback;
            crc[16]      = crc[17];
            crc[17]      = crc[18];
            crc[18]      = crc[19];
            crc[19]      = crc[20] ^ crc_feedback;
            crc[20]      = crc[21] ^ crc_feedback;
            crc[21]      = crc[22] ^ crc_feedback;
            crc[22]      = crc[23];
            crc[23]      = crc[24] ^ crc_feedback;
            crc[24]      = crc[25] ^ crc_feedback;
            crc[25]      = crc[26];
            crc[26]      = crc[27] ^ crc_feedback;
            crc[27]      = crc[28] ^ crc_feedback;
            crc[28]      = crc[29];
            crc[29]      = crc[30] ^ crc_feedback;
            crc[30]      = crc[31] ^ crc_feedback;
            crc[31]      =           crc_feedback;
        end

        // return the CRC result
        fcs = ~ crc;

    end
    endtask // calc_crc

    //----------------------------------------------------------------------------
    // Test Bench signals and constanggs
    //----------------------------------------------------------------------------

    // Delay to provide setup and hold timing at the GMII/RGMII.
    parameter dly = 2;  // 2 ns

    parameter gtx_period = 10;  // ns

    parameter SEQ_OFFSET = 14;


    // testbench signals
    
    wire        gtx_clk;
    reg         mmcm_clk_in;
    reg         reset;
    reg  [3:0]  demo_mode_error = 1'b0;

    wire [3:0]  mdc;
    wire [3:0]  mdio;
    reg  [5:0]  mdio_count [0:3];
    reg  [3:0]  last_mdio;
    reg  [3:0]  mdio_read;
    reg  [3:0]  mdio_addr;
    reg  [3:0]  mdio_fail;
    wire [3:0]  rgmii_txc;
    wire [3:0]  rgmii_tx_ctl;
    wire [3:0]  rgmii_txd [0:3];
    reg  [3:0]  rgmii_rxc_1000;
    reg  [3:0]  rgmii_rxc_100;
    reg  [3:0]  rgmii_rxc_10;
    wire [3:0]  rgmii_rxc;
    reg  [3:0]  rgmii_rx_ctl;
    reg  [3:0]  rgmii_rxd [0:3];
    wire [3:0]  inband_link_status;
    wire [1:0]  inband_clock_speed [0:3];
    wire [3:0]  inband_duplex_status;

    // testbench control semaphores
    reg         rx_stimulus_warmup_finished;
    reg [3:0]   rx_stimulus_pressure_finished;
    reg [3:0]   tx_monitor_finished_1G;
    reg [3:0]   tx_monitor_finished_10M;
    reg [3:0]   tx_monitor_finished_100M;
    reg [3:0]   management_config_finished;

    reg [1:0]   phy_speed [0:3];
    reg [1:0]   mac_speed [0:3];
    reg [3:0]   update_speed;

    wire [3:0]  rgmii_rx_ctl_dut;
    wire [3:0]  rgmii_rxd_dut [0:3];

    reg [3:0]   gen_tx_data;
    reg [3:0]   check_tx_data;
    reg [3:0]   config_bist;
    
    wire [3:0]  frame_error;
    reg  [3:0]  bist_mode_error;
    wire [3:0]  serial_response;

    reg [3:0]   count_frame;
    reg [3:0]   vlan_frame [0:3] ;
    reg [16:0]  vlan_count [0:3];
    reg [16:0]  total_count [0:3];

    // Generate a delayed rgmii_rxc to match the spec
    wire [3:0]  delay_rxc;
    wire [3:0]  delay_rxc_lcl;
    assign #2 delay_rxc_lcl = rgmii_rxc;
    // only want the delay if the rgmii isn't looped back
    // assign       delay_rxc = (TB_MODE == "BIST") ? rgmii_txc : delay_rxc_lcl;
    assign delay_rxc = delay_rxc_lcl;

    // select between loopback or local data
    // assign rgmii_rxd_dut    = (TB_MODE == "BIST") ? rgmii_txd    : rgmii_rxd;
    // assign rgmii_rx_ctl_dut = (TB_MODE == "BIST") ? rgmii_tx_ctl : rgmii_rx_ctl;
    // assign rgmii_rxd_dut = rgmii_rxd;
    // assign rgmii_rx_ctl_dut = rgmii_rx_ctl;

    //----------------------------------------------------------------------------
    // Wire up Device Under Test
    //----------------------------------------------------------------------------

    tns_tsn_03 dut (
        .glbl_rstn                  (!reset),
        .sys_clk                    (mmcm_clk_in),
//        .gtx_clk_bufg_out           (gtx_clk),
        .rgmii_txd_flat             ({rgmii_txd[3], rgmii_txd[2], rgmii_txd[1], rgmii_txd[0]}),
        .rgmii_tx_ctl               (rgmii_tx_ctl),
        .rgmii_txc                  (rgmii_txc),
        .rgmii_rxd_flat             ({rgmii_rxd[3], rgmii_rxd[2], rgmii_rxd[1], rgmii_rxd[0]}),
        .rgmii_rx_ctl               (rgmii_rx_ctl),
        .rgmii_rxc                  (delay_rxc),
        .mdio                       (mdio),
        .mdc                        (mdc)
    );


    //---------------------------------------------------------------------------
    //-- If the simulation is still going then
    //-- something has gone wrong
    //---------------------------------------------------------------------------
    //    initial
    //    begin
    //        #680000000;
    //        $display("** ERROR: Simulation Running Forever");
    //        $stop;
    //    end

    //----------------------------------------------------------------------------
    // Simulate the MDIO -
    // respond with sensible data to mdio reads and accept writes
    //----------------------------------------------------------------------------
    // expect mdio to try and read from reg addr 1 - return all 1's if we don't
    // want any other mdio accesses
    // if any other response then mdio will write to reg_addr 9 then 4 then 0
    // (may check for expected write data?)
    // finally mdio read from reg addr 1 until bit 5 is seen high
    // NOTE - do not check any other bits so could drive all high again..


    // count through the mdio transfer
    genvar i;
    generate
        for (i = 0; i < 4; i = i + 1)
        begin
            always @(posedge mdc[i] or posedge reset)
            begin
                if (reset) begin
                    mdio_count[i] <= 0;
                    last_mdio[i] <= 1'b0;
                end
                else begin
                    last_mdio[i] <= mdio[i];
                    if (mdio_count[i] >= 32) begin
                    mdio_count[i] <= 0;
                    end
                    else if (mdio_count[i] != 0) begin
                    mdio_count[i] <= mdio_count[i] + 1;
                    end
                    else begin // only get here if mdio state is 0 - now look for a start
                    if ((mdio[i] === 1'b1) && (last_mdio[i] === 1'b0))
                        mdio_count[i] <= 1;
                    end
                end
            end
            assign mdio[i] = (mdio_read[i] & (mdio_count[i] >= 14) & (mdio_count[i] <= 31)) ? 1'b1 : 1'bz;

            // only respond to phy addr 7 and reg address == 1 (PHY_STATUS)
            always @(posedge mdc[i] or posedge reset)
            begin
                if (reset) begin
                    mdio_read[i] <= 1'b0;
                    mdio_addr[i] <= 1'b1; // this will go low if the address doesn't match required
                    mdio_fail[i] <= 1'b0;
                end
                else
                begin
                    if (mdio_count[i] == 2) begin
                    mdio_addr[i] <= 1'b1;    // new access so address needs to be revalidated
                    if ({last_mdio[i],mdio[i]} === 2'b10)
                        mdio_read[i] <= 1'b1;
                    else // take a write as a default as won't drive at the wrong time
                        mdio_read[i] <= 1'b0;
                    end
                    else if ((mdio_count[i] <= 12)) begin
                    // check address is phy addr/reg addr are correct
                    if (mdio_count[i] <= 7 & mdio_count[i] >= 5) begin
                        if (mdio[i] !== 1'b1)
                            mdio_addr[i] <= 1'b0;
                    end
                    else begin
                        if (mdio[i] !== 1'b0)
                            mdio_addr[i] <= 1'b0;
                    end
                    end
                    else if ((mdio_count[i] == 14)) begin
                    if (!mdio_read[i] & (mdio[i] | !last_mdio[i])) begin
                        $display("FAIL : Write TA phase is incorrect at %t ps", $time);
                    end
                    end
                    else if ((mdio_count[i] >= 15) & (mdio_count[i] <= 30) & mdio_addr[i]) begin
                    if (!mdio_read[i]) begin
                        if (mdio_count[i] == 20) begin
                            if (mdio[i]) begin
                                mdio_fail[i] <= 1;
                                $display("FAIL : Expected bit 10 of mdio write data to be 0 at %t ps", $time);
                            end
                        end
                        else begin
                            if (!mdio[i]) begin
                                mdio_fail[i] <= 1;
                                $display("FAIL : Expected all except bit 10 of mdio write data to be 1 at %t ps", $time);
                            end
                        end
                    end
                    end
                end
            end
        end
    endgenerate


    //----------------------------------------------------------------------------
    // Clock drivers
    //----------------------------------------------------------------------------
    

    //drives input to an MMCM at 50MHz which creates gtx_clk at 125 MHz
    initial
    begin
        
        mmcm_clk_in <= 1'b0;
        
    #80;
        forever
        begin
        mmcm_clk_in <= 1'b0;
        
        #gtx_period;
        mmcm_clk_in <= 1'b1;
        
        #gtx_period;
        end
    end

        

    // drives rgmii_rxc_1000 at 125 MHz
    initial
    begin
        rgmii_rxc_1000 <= 4'b0000;
        #10;
        forever
        begin
        rgmii_rxc_1000 <= 4'b0000;
        #4;
        rgmii_rxc_1000 <= 4'b1111;
        #4;
        end
    end


    // drives rgmii_rxc_100 at 25 MHz
    initial
    begin
        rgmii_rxc_100 <= 4'b0000;
        #10;
        forever
        begin
        rgmii_rxc_100 <= 4'b0000;
        #20;
        rgmii_rxc_100 <= 4'b1111;
        #20;
        end
    end


    // drives rgmii_rxc_10 at 2.5 MHz
    initial
    begin
        rgmii_rxc_10 <= 4'b0000;
        #10;
        forever
        begin
        rgmii_rxc_10 <= 4'b0000;
        #200;
        rgmii_rxc_10 <= 4'b1111;
        #200;
        end
    end

    // want a clean swicth between the clocks - provide a low setting
    // Select between 10Mb/s, 100Mb/s and 1Gb/s RGMII Rx clock frequencies
    assign rgmii_rxc[0] = (phy_speed[0] == 2'b11 ? 1'b0 :
                        phy_speed[0] == 2'b10 ? rgmii_rxc_1000[0] :
                        (phy_speed[0] == 2'b01 ? rgmii_rxc_100[0] : rgmii_rxc_10[0]));
    assign rgmii_rxc[1] = (phy_speed[1] == 2'b11 ? 1'b0 :
                        phy_speed[1] == 2'b10 ? rgmii_rxc_1000[1] :
                        (phy_speed[1] == 2'b01 ? rgmii_rxc_100[1] : rgmii_rxc_10[1]));
    assign rgmii_rxc[2] = (phy_speed[2] == 2'b11 ? 1'b0 :
                        phy_speed[2] == 2'b10 ? rgmii_rxc_1000[2] :
                        (phy_speed[2] == 2'b01 ? rgmii_rxc_100[2] : rgmii_rxc_10[2]));
    assign rgmii_rxc[3] = (phy_speed[3] == 2'b11 ? 1'b0 :
                        phy_speed[3] == 2'b10 ? rgmii_rxc_1000[3] :
                        (phy_speed[3] == 2'b01 ? rgmii_rxc_100[3] : rgmii_rxc_10[3]));

    //----------------------------------------------------------------------------
    // A Task to reset the MAC
    //----------------------------------------------------------------------------
    task mac_reset;
        begin
        $display("** Note: Resetting core...");

        reset <= 1'b1;
        #400

        reset <= 1'b0;

        $display("** Note: Timing checks are valid");
        end
    endtask // mac_reset;
    
    generate
        for (i = 0; i < 4; i = i + 1)
        begin
            // count vlan frame bytes
            always @(posedge gtx_clk or posedge reset)
            begin
                if (reset) begin
                    count_frame[i] <= 0;
                end
                else if (vlan_frame[i])
                    count_frame[i] <= 1;
                else if (!rgmii_tx_ctl[i])
                    count_frame[i] <= 0;
            end

            // count vlan frame bytes
            always @(posedge gtx_clk or posedge reset)
            begin
                if (reset) begin
                    vlan_count[i] <= 0;
                end
                else if (vlan_frame[i])
                    vlan_count[i] <= vlan_count[i] + 12 + 8 + 12; // only detect vlan frame after 12 bytes - also aloow for preamble and ifg
                else if (count_frame[i])
                    vlan_count[i] <= vlan_count[i] + 1;
            end

            // count possible frame bytes - only start when first vlan frame seen (avoids reset gap)
            always @(posedge gtx_clk or posedge reset)
            begin
                if (reset) begin
                    total_count[i] <= 0;
                end
                else if (|total_count[i])
                    total_count[i] <= total_count[i] + 1;
                else if (vlan_frame[i])
                    total_count[i] <= total_count[i] + 12 + 8 + 12;
            end

            // monitor frame error and output error when asserted (with timestamp)
            always @(posedge gtx_clk or posedge reset)
            begin
                if (reset) begin
                    bist_mode_error[i] <= 0;
                end
                    
                else if (frame_error[i] & !bist_mode_error[i]) begin
                    bist_mode_error[i] <= 1;
                    $display("ERROR: frame mismatch at time %t ps", $time);
                end
            end
            
        end
    endgenerate


    //----------------------------------------------------------------------------
    // Management process. This process waits for setup to complete by monitoring the mdio
    // (the host always runs at gtx_clk so the setup after mdio accesses are complete
    // doesn't take long) and then allows packets to be sent
    //----------------------------------------------------------------------------
    
    reg [3:0] wait_mdio_count_32 = 4'b0;
    reg [3:0] wait_mdio_count_0 = 4'b0;
    
    initial
    begin : p_management

        mac_speed[0] <= 2'b01;
        mac_speed[1] <= 2'b01;
        mac_speed[2] <= 2'b01;
        mac_speed[3] <= 2'b01;
                        
        phy_speed[0] <= 2'b01;
        phy_speed[1] <= 2'b01;
        phy_speed[2] <= 2'b01;
        phy_speed[3] <= 2'b01;

        update_speed <= 4'b0;
        gen_tx_data <= 4'b0;
        check_tx_data <= 4'b0;
        config_bist <= 4'b0;
        management_config_finished <= 4'b0;

        // reset the core
        mac_reset;


        // check mdio
        // wait for the mdio access and remainder of setup accesses (internal)
        while (wait_mdio_count_0[2:0] !== 3'b111)
        begin
            @(mdio_count[0] or mdio_count[1] or mdio_count[2] or mdio_count[3]) begin
                if (mdio_count[0] == 32) begin
                    wait_mdio_count_32[0] = 1;
                end
                if (mdio_count[1] == 32) begin
                    wait_mdio_count_32[1] = 1;
                end
                if (mdio_count[2] == 32) begin
                    wait_mdio_count_32[2] = 1;
                end
                if (mdio_count[3] == 32) begin
                    wait_mdio_count_32[3] = 1;
                end
                if ((mdio_count[0] == 0) && (wait_mdio_count_32[0] == 1)) begin
                    wait_mdio_count_0[0] = 1;
                end
                if ((mdio_count[1] == 0) && (wait_mdio_count_32[1] == 1)) begin
                    wait_mdio_count_0[1] = 1;
                end
                if ((mdio_count[2] == 0) && (wait_mdio_count_32[2] == 1)) begin
                    wait_mdio_count_0[2] = 1;
                end
                if ((mdio_count[3] == 0) && (wait_mdio_count_32[3] == 1)) begin
                    wait_mdio_count_0[3] = 1;
                end
            end
        end

        // wait (mdio_count == 32);
        // wait (mdio_count == 0);

        // Signal that configuration is complete.  Other processes will now
        // be allowed to run.
        management_config_finished = 4'b1111;

        // The stimulus process will now send 5 frames at 1Gb/s.
        //------------------------------------------------------------------

        // Wait for 1G monitor process to complete.
        // wait (tx_monitor_finished_1G == 4'b1111);
        wait (rx_stimulus_pressure_finished == 4'b1111);
        // #100000000
        

        // Our work here is done
        // if (demo_mode_error == 4'b0 && bist_mode_error == 4'b0) begin
        //     $display("Test completed successfully");
        // end
        // $display("Simulation Stopped");
        // $stop;
    end // p_management



    //----------------------------------------------------------------------------
    // Procedure to inject a frame into the receiver at 1Gb/s
    //----------------------------------------------------------------------------
    task automatic send_frame_1g_port0;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_0.frombits(frame);
        rx_stimulus_working_frame_0.data[SEQ_OFFSET] = seq_num[31:24];
        rx_stimulus_working_frame_0.data[SEQ_OFFSET + 1] = seq_num[23:16];
        rx_stimulus_working_frame_0.data[SEQ_OFFSET + 2] = seq_num[15:8];
        rx_stimulus_working_frame_0.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[0]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[0]   <= 4'h5;
            rgmii_rx_ctl[0] <= 1'b1;
            @(rgmii_rxc[0]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[0] <= 4'h5;
        rgmii_rx_ctl[0] <= 1'b1;
        @(rgmii_rxc[0])
        rgmii_rxd[0] <= 4'hD;
        rgmii_rx_ctl[0] <= 1'b1;
        @(rgmii_rxc[0])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_0.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[0]    <= rx_stimulus_working_frame_0.data[column_index][3:0];
            rgmii_rx_ctl[0] <= rx_stimulus_working_frame_0.valid[column_index];
            @(rgmii_rxc[0])
            rgmii_rxd[0]    <= rx_stimulus_working_frame_0.data[column_index][7:4];
            rgmii_rx_ctl[0] <= rx_stimulus_working_frame_0.valid[column_index] ^ rx_stimulus_working_frame_0.error[column_index];
            calc_crc(rx_stimulus_working_frame_0.data[column_index], fcs);

            column_index = column_index + 1;
            @(rgmii_rxc[0]);  // wait for next clock tick

        end

        $display("port0 send %d bytes.", column_index);

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[0]    <= fcs[3:0];
            1 : rgmii_rxd[0]    <= fcs[11:8];
            2 : rgmii_rxd[0]    <= fcs[19:16];
            3 : rgmii_rxd[0]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[0] <= 1'b1;
            @(rgmii_rxc[0])
            case(I)
            0 : rgmii_rxd[0]    <= fcs[7:4];
            1 : rgmii_rxd[0]    <= fcs[15:12];
            2 : rgmii_rxd[0]    <= fcs[23:20];
            3 : rgmii_rxd[0]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[0] <= 1'b1;

            @(rgmii_rxc[0]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[0]       <= 4'h0;
        rgmii_rx_ctl[0]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        // TODO on wiki, it is 12 octets.
        for (I = 0; I < 16; I = I + 1)
            @(rgmii_rxc[0]);
        // $display("send one frame from port 0, 1g, CRC %h.", fcs);

        // for (I = 0; I < 27000; I = I + 1)
        //     @(rgmii_rxc[0]);

        end
        
        
    endtask // send_frame_1g;

    task automatic send_frame_1g_port1;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_1.frombits(frame);

        rx_stimulus_working_frame_1.data[SEQ_OFFSET] = seq_num[31:24];
        rx_stimulus_working_frame_1.data[SEQ_OFFSET + 1] = seq_num[23:16];
        rx_stimulus_working_frame_1.data[SEQ_OFFSET + 2] = seq_num[15:8];
        rx_stimulus_working_frame_1.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[1]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[1]   <= 4'h5;
            rgmii_rx_ctl[1] <= 1'b1;
            @(rgmii_rxc[1]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[1] <= 4'h5;
        rgmii_rx_ctl[1] <= 1'b1;
        @(rgmii_rxc[1])
        rgmii_rxd[1] <= 4'hD;
        rgmii_rx_ctl[1] <= 1'b1;
        @(rgmii_rxc[1])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_1.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[1]    <= rx_stimulus_working_frame_1.data[column_index][3:0];
            rgmii_rx_ctl[1] <= rx_stimulus_working_frame_1.valid[column_index];
            @(rgmii_rxc[1])
            rgmii_rxd[1]    <= rx_stimulus_working_frame_1.data[column_index][7:4];
            rgmii_rx_ctl[1] <= rx_stimulus_working_frame_1.valid[column_index] ^ rx_stimulus_working_frame_1.error[column_index];
            calc_crc(rx_stimulus_working_frame_1.data[column_index], fcs);

            column_index = column_index + 1;
            @(rgmii_rxc[1]);  // wait for next clock tick

        end

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[1]    <= fcs[3:0];
            1 : rgmii_rxd[1]    <= fcs[11:8];
            2 : rgmii_rxd[1]    <= fcs[19:16];
            3 : rgmii_rxd[1]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[1] <= 1'b1;
            @(rgmii_rxc[1])
            case(I)
            0 : rgmii_rxd[1]    <= fcs[7:4];
            1 : rgmii_rxd[1]    <= fcs[15:12];
            2 : rgmii_rxd[1]    <= fcs[23:20];
            3 : rgmii_rxd[1]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[1] <= 1'b1;

            @(rgmii_rxc[1]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[1]       <= 4'h0;
        rgmii_rx_ctl[1]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        for (I = 0; I < 16; I = I + 1)
            @(rgmii_rxc[1]);
        // for (I = 0; I < 27000; I = I + 1)
        //     @(rgmii_rxc[1]);

        end
    endtask // send_frame_1g;

    task automatic send_frame_1g_port2;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_2.frombits(frame);
        rx_stimulus_working_frame_2.data[SEQ_OFFSET] = seq_num[31:24];
        rx_stimulus_working_frame_2.data[SEQ_OFFSET + 1] = seq_num[23:16];
        rx_stimulus_working_frame_2.data[SEQ_OFFSET + 2] = seq_num[15:8];
        rx_stimulus_working_frame_2.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[2]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[2]   <= 4'h5;
            rgmii_rx_ctl[2] <= 1'b1;
            @(rgmii_rxc[2]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[2] <= 4'h5;
        rgmii_rx_ctl[2] <= 1'b1;
        @(rgmii_rxc[2])
        rgmii_rxd[2] <= 4'hD;
        rgmii_rx_ctl[2] <= 1'b1;
        @(rgmii_rxc[2])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_2.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[2]    <= rx_stimulus_working_frame_2.data[column_index][3:0];
            rgmii_rx_ctl[2] <= rx_stimulus_working_frame_2.valid[column_index];
            @(rgmii_rxc[2])
            rgmii_rxd[2]    <= rx_stimulus_working_frame_2.data[column_index][7:4];
            rgmii_rx_ctl[2] <= rx_stimulus_working_frame_2.valid[column_index] ^ rx_stimulus_working_frame_2.error[column_index];
            calc_crc(rx_stimulus_working_frame_2.data[column_index], fcs);

            column_index = column_index + 1;
            @(rgmii_rxc[2]);  // wait for next clock tick

        end

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[2]    <= fcs[3:0];
            1 : rgmii_rxd[2]    <= fcs[11:8];
            2 : rgmii_rxd[2]    <= fcs[19:16];
            3 : rgmii_rxd[2]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[2] <= 1'b1;
            @(rgmii_rxc[2])
            case(I)
            0 : rgmii_rxd[2]    <= fcs[7:4];
            1 : rgmii_rxd[2]    <= fcs[15:12];
            2 : rgmii_rxd[2]    <= fcs[23:20];
            3 : rgmii_rxd[2]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[2] <= 1'b1;

            @(rgmii_rxc[2]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[2]       <= 4'h0;
        rgmii_rx_ctl[2]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        for (I = 0; I < 16; I = I + 1)
            @(rgmii_rxc[2]);
        // for (I = 0; I < 27000; I = I + 1)
        //     @(rgmii_rxc[2]);

        end
    endtask // send_frame_1g;

    task automatic send_frame_1g_port3;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_3.frombits(frame);
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET] = seq_num[31:24];
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET + 1] = seq_num[23:16];
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET + 2] = seq_num[15:8];
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[3]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[3]   <= 4'h5;
            rgmii_rx_ctl[3] <= 1'b1;
            @(rgmii_rxc[3]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[3] <= 4'h5;
        rgmii_rx_ctl[3] <= 1'b1;
        @(rgmii_rxc[3])
        rgmii_rxd[3] <= 4'hD;
        rgmii_rx_ctl[3] <= 1'b1;
        @(rgmii_rxc[3])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_3.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[3]    <= rx_stimulus_working_frame_3.data[column_index][3:0];
            rgmii_rx_ctl[3] <= rx_stimulus_working_frame_3.valid[column_index];
            @(rgmii_rxc[3])
            rgmii_rxd[3]    <= rx_stimulus_working_frame_3.data[column_index][7:4];
            rgmii_rx_ctl[3] <= rx_stimulus_working_frame_3.valid[column_index] ^ rx_stimulus_working_frame_3.error[column_index];
            calc_crc(rx_stimulus_working_frame_3.data[column_index], fcs);

            column_index = column_index + 1;
            @(rgmii_rxc[3]);  // wait for next clock tick

        end

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[3]    <= fcs[3:0];
            1 : rgmii_rxd[3]    <= fcs[11:8];
            2 : rgmii_rxd[3]    <= fcs[19:16];
            3 : rgmii_rxd[3]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[3] <= 1'b1;
            @(rgmii_rxc[3])
            case(I)
            0 : rgmii_rxd[3]    <= fcs[7:4];
            1 : rgmii_rxd[3]    <= fcs[15:12];
            2 : rgmii_rxd[3]    <= fcs[23:20];
            3 : rgmii_rxd[3]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[3] <= 1'b1;

            @(rgmii_rxc[3]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[3]       <= 4'h0;
        rgmii_rx_ctl[3]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        for (I = 0; I < 16; I = I + 1)
            @(rgmii_rxc[3]);
        // for (I = 0; I < 27000; I = I + 1)
        //     @(rgmii_rxc[3]);

        end
    endtask // send_frame_1g;


    //----------------------------------------------------------------------------
    // Procedure to inject a frame into the receiver at 100Mb/s
    //----------------------------------------------------------------------------
    task automatic send_frame_100m_port0;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_0.frombits(frame);
        rx_stimulus_working_frame_0.data[SEQ_OFFSET] = seq_num[31:24];
        rx_stimulus_working_frame_0.data[SEQ_OFFSET + 1] = seq_num[23:16];
        rx_stimulus_working_frame_0.data[SEQ_OFFSET + 2] = seq_num[15:8];
        rx_stimulus_working_frame_0.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[0]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[0]   <= 4'h5;
            rgmii_rx_ctl[0] <= 1'b1;
            @(posedge rgmii_rxc[0]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[0] <= 4'h5;
        rgmii_rx_ctl[0] <= 1'b1;
        @(posedge rgmii_rxc[0]);
        rgmii_rxd[0] <= 4'hD;
        rgmii_rx_ctl[0] <= 1'b1;
        @(posedge rgmii_rxc[0]);

        // loop over columns in frame.
        while (rx_stimulus_working_frame_0.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[0]    <= rx_stimulus_working_frame_0.data[column_index][3:0];
            rgmii_rx_ctl[0] <= rx_stimulus_working_frame_0.valid[column_index];
            @(posedge rgmii_rxc[0])
            rgmii_rxd[0]    <= rx_stimulus_working_frame_0.data[column_index][7:4];
            rgmii_rx_ctl[0] <= rx_stimulus_working_frame_0.valid[column_index] ^ rx_stimulus_working_frame_0.error[column_index];
            calc_crc(rx_stimulus_working_frame_0.data[column_index], fcs);

            column_index = column_index + 1;
            @(posedge rgmii_rxc[0]);  // wait for next clock tick

        end

        $display("port0 send %d bytes.", column_index);

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[0]    <= fcs[3:0];
            1 : rgmii_rxd[0]    <= fcs[11:8];
            2 : rgmii_rxd[0]    <= fcs[19:16];
            3 : rgmii_rxd[0]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[0] <= 1'b1;
            @(posedge rgmii_rxc[0])
            case(I)
            0 : rgmii_rxd[0]    <= fcs[7:4];
            1 : rgmii_rxd[0]    <= fcs[15:12];
            2 : rgmii_rxd[0]    <= fcs[23:20];
            3 : rgmii_rxd[0]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[0] <= 1'b1;

            @(posedge rgmii_rxc[0]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[0]       <= 4'h0;
        rgmii_rx_ctl[0]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        // TODO on wiki, it is 12 octets.
        for (I = 0; I < 32; I = I + 1)
            @(rgmii_rxc[0]);
        // $display("send one frame from port 0, 1g, CRC %h.", fcs);

    

        end
        
        
    endtask // send_frame_1g;

    task automatic send_frame_100m_port1;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_1.frombits(frame);

        rx_stimulus_working_frame_1.data[SEQ_OFFSET] = seq_num[31:24];
        rx_stimulus_working_frame_1.data[SEQ_OFFSET + 1] = seq_num[23:16];
        rx_stimulus_working_frame_1.data[SEQ_OFFSET + 2] = seq_num[15:8];
        rx_stimulus_working_frame_1.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[1]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[1]   <= 4'h5;
            rgmii_rx_ctl[1] <= 1'b1;
            @(posedge rgmii_rxc[1]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[1] <= 4'h5;
        rgmii_rx_ctl[1] <= 1'b1;
        @(posedge rgmii_rxc[1])
        rgmii_rxd[1] <= 4'hD;
        rgmii_rx_ctl[1] <= 1'b1;
        @(posedge rgmii_rxc[1])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_1.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[1]    <= rx_stimulus_working_frame_1.data[column_index][3:0];
            rgmii_rx_ctl[1] <= rx_stimulus_working_frame_1.valid[column_index];
            @(posedge rgmii_rxc[1])
            rgmii_rxd[1]    <= rx_stimulus_working_frame_1.data[column_index][7:4];
            rgmii_rx_ctl[1] <= rx_stimulus_working_frame_1.valid[column_index] ^ rx_stimulus_working_frame_1.error[column_index];
            calc_crc(rx_stimulus_working_frame_1.data[column_index], fcs);

            column_index = column_index + 1;
            @(posedge rgmii_rxc[1]);  // wait for next clock tick

        end

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[1]    <= fcs[3:0];
            1 : rgmii_rxd[1]    <= fcs[11:8];
            2 : rgmii_rxd[1]    <= fcs[19:16];
            3 : rgmii_rxd[1]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[1] <= 1'b1;
            @(posedge rgmii_rxc[1])
            case(I)
            0 : rgmii_rxd[1]    <= fcs[7:4];
            1 : rgmii_rxd[1]    <= fcs[15:12];
            2 : rgmii_rxd[1]    <= fcs[23:20];
            3 : rgmii_rxd[1]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[1] <= 1'b1;

            @(posedge rgmii_rxc[1]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[1]       <= 4'h0;
        rgmii_rx_ctl[1]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        for (I = 0; I < 32; I = I + 1)
            @(rgmii_rxc[1]);

        end
    endtask // send_frame_100m_port1;

    task automatic send_frame_100m_port2;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_2.frombits(frame);
        rx_stimulus_working_frame_2.data[SEQ_OFFSET] = seq_num[31:24];
        rx_stimulus_working_frame_2.data[SEQ_OFFSET + 1] = seq_num[23:16];
        rx_stimulus_working_frame_2.data[SEQ_OFFSET + 2] = seq_num[15:8];
        rx_stimulus_working_frame_2.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[2]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[2]   <= 4'h5;
            rgmii_rx_ctl[2] <= 1'b1;
            @(posedge rgmii_rxc[2]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[2] <= 4'h5;
        rgmii_rx_ctl[2] <= 1'b1;
        @(posedge rgmii_rxc[2])
        rgmii_rxd[2] <= 4'hD;
        rgmii_rx_ctl[2] <= 1'b1;
        @(posedge rgmii_rxc[2])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_2.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[2]    <= rx_stimulus_working_frame_2.data[column_index][3:0];
            rgmii_rx_ctl[2] <= rx_stimulus_working_frame_2.valid[column_index];
            @(posedge rgmii_rxc[2])
            rgmii_rxd[2]    <= rx_stimulus_working_frame_2.data[column_index][7:4];
            rgmii_rx_ctl[2] <= rx_stimulus_working_frame_2.valid[column_index] ^ rx_stimulus_working_frame_2.error[column_index];
            calc_crc(rx_stimulus_working_frame_2.data[column_index], fcs);

            column_index = column_index + 1;
            @(posedge rgmii_rxc[2]);  // wait for next clock tick

        end

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[2]    <= fcs[3:0];
            1 : rgmii_rxd[2]    <= fcs[11:8];
            2 : rgmii_rxd[2]    <= fcs[19:16];
            3 : rgmii_rxd[2]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[2] <= 1'b1;
            @(posedge rgmii_rxc[2])
            case(I)
            0 : rgmii_rxd[2]    <= fcs[7:4];
            1 : rgmii_rxd[2]    <= fcs[15:12];
            2 : rgmii_rxd[2]    <= fcs[23:20];
            3 : rgmii_rxd[2]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[2] <= 1'b1;

            @(posedge rgmii_rxc[2]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[2]       <= 4'h0;
        rgmii_rx_ctl[2]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        for (I = 0; I < 32; I = I + 1)
            @(rgmii_rxc[2]);

        end
    endtask // send_frame_100m_port2;

    task automatic send_frame_100m_port3;
        input   `FRAME_TYP frame;
        input integer seq_num;
        integer column_index;
        integer I;
        reg [31:0] fcs;
        begin
        // import the frame into scratch space
        rx_stimulus_working_frame_3.frombits(frame);
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET] = seq_num[31:24];
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET + 1] = seq_num[23:16];
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET + 2] = seq_num[15:8];
        // rx_stimulus_working_frame_3.data[SEQ_OFFSET + 3] = seq_num[7:0];

        // Reset the FCS calculation
        fcs = 32'b0;
        @(posedge rgmii_rxc[3]);

        column_index = 0;

        // Adding the preamble field
        for (I = 0; I <= 13; I = I + 1)
        begin
            rgmii_rxd[3]   <= 4'h5;
            rgmii_rx_ctl[3] <= 1'b1;
            @(posedge rgmii_rxc[3]);
        end

        // Adding the Start of Frame Delimiter (SFD)
        rgmii_rxd[3] <= 4'h5;
        rgmii_rx_ctl[3] <= 1'b1;
        @(posedge rgmii_rxc[3])
        rgmii_rxd[3] <= 4'hD;
        rgmii_rx_ctl[3] <= 1'b1;
        @(posedge rgmii_rxc[3])

        // loop over columns in frame.
        while (rx_stimulus_working_frame_3.valid[column_index] !== 1'b0)
        begin
            // send one column of data
            rgmii_rxd[3]    <= rx_stimulus_working_frame_3.data[column_index][3:0];
            rgmii_rx_ctl[3] <= rx_stimulus_working_frame_3.valid[column_index];
            @(posedge rgmii_rxc[3])
            rgmii_rxd[3]    <= rx_stimulus_working_frame_3.data[column_index][7:4];
            rgmii_rx_ctl[3] <= rx_stimulus_working_frame_3.valid[column_index] ^ rx_stimulus_working_frame_3.error[column_index];
            calc_crc(rx_stimulus_working_frame_3.data[column_index], fcs);

            column_index = column_index + 1;
            @(posedge rgmii_rxc[3]);  // wait for next clock tick

        end

        // Send the CRC.
        for (I = 0; I < 4; I = I + 1)
        begin
            case(I)
            0 : rgmii_rxd[3]    <= fcs[3:0];
            1 : rgmii_rxd[3]    <= fcs[11:8];
            2 : rgmii_rxd[3]    <= fcs[19:16];
            3 : rgmii_rxd[3]    <= fcs[27:24];
            endcase
            rgmii_rx_ctl[3] <= 1'b1;
            @(posedge rgmii_rxc[3])
            case(I)
            0 : rgmii_rxd[3]    <= fcs[7:4];
            1 : rgmii_rxd[3]    <= fcs[15:12];
            2 : rgmii_rxd[3]    <= fcs[23:20];
            3 : rgmii_rxd[3]    <= fcs[31:28];
            endcase
            rgmii_rx_ctl[3] <= 1'b1;

            @(posedge rgmii_rxc[3]);  // wait for next clock tick
        end

        // Clear the data lines.
        rgmii_rxd[3]       <= 4'h0;
        rgmii_rx_ctl[3]    <= 1'b0;

        // Adding the minimum Interframe gap for a receiver (8 idles)
        for (I = 0; I < 32; I = I + 1)
            @(rgmii_rxc[3]);

        end
    endtask // send_frame_100m_port3;




    // Stimulus process: warm up.
    initial 
    begin: p_rx_stimulus_warmup
        rx_stimulus_warmup_finished = 0;
        rx_stimulus_pressure_finished = 4'b0;

        rgmii_rxd[0]      = 4'h0;
        rgmii_rxd[1]      = 4'h0;
        rgmii_rxd[2]      = 4'h0;
        rgmii_rxd[3]      = 4'h0;

        rgmii_rx_ctl   = 4'b0000;
        
        while (management_config_finished !== 4'hf)
        // wait for the internal resets to settle before staring to send traffic
        #800;
        // $display("Rx Stimulus warm up.");
        // if (mac_speed[0] == 2'b10) begin
        //     send_frame_1g_port0(frame0.tobits(0), -1);
        // end
        // else if(mac_speed[0] == 2'b01) begin
        //     send_frame_100m_port0(frame0.tobits(0), -1);
        // end
        // #10;
        // if (mac_speed[1] == 2'b10) begin
        //     send_frame_1g_port1(frame2.tobits(0), -1);
        // end
        // else if(mac_speed[1] == 2'b01) begin
        //     send_frame_100m_port1(frame2.tobits(0), -1);
        // end
        // #10;
        // if (mac_speed[2] == 2'b10) begin
        //     send_frame_1g_port2(frame3.tobits(0), -1);
        // end
        // else if(mac_speed[2] == 2'b01) begin
        //     send_frame_100m_port2(frame3.tobits(0), -1);
        // end
        // #10;
        // if (mac_speed[3] == 2'b10) begin
        //     send_frame_1g_port3(frame1.tobits(0), -1);
        // end
        // else if(mac_speed[3] == 2'b01) begin
        //     send_frame_100m_port3(frame1.tobits(0), -1);
        // end
        // #10;
        // $display("Warmup done.");
        rx_stimulus_warmup_finished = 1;
        // wait (tx_monitor_finished_1G == 4'b1111);
    end

    integer i_stimulus_port0;

    initial
    begin : p_rx_stimulus_port0
        wait(rx_stimulus_warmup_finished == 1);
        #10;

        // 1 Gb/s speed
        //-----------------------------------------------------
        
        // Presure test
        // $display("Phase two of stimulation port 0: Noting, just receive.");
        for (i_stimulus_port0 = 0; i_stimulus_port0 < 100; i_stimulus_port0 = i_stimulus_port0 + 1) begin
            $display ("Port 0 Send: 1->4 #0d", i_stimulus_port0);
            if (mac_speed[0] == 2'b10) begin
                send_frame_1g_port0(frame0.tobits(0), i_stimulus_port0);
            end
            else if (mac_speed[0] == 2'b01) begin
                send_frame_100m_port0(frame0.tobits(0), i_stimulus_port0);
            end
        end

        // wait (tx_monitor_finished_1G == 4'b1111);
        rx_stimulus_pressure_finished[0] = 1;
        #10;
    end // p_rx_stimulus_port0

    integer i_stimulus_port1;

    initial
    begin : p_rx_stimulus_port1
        wait(rx_stimulus_warmup_finished == 1);
        #10;

        // 1 Gb/s speed
        //-----------------------------------------------------
        
        // Presure test
        $display("Phase two of stimulation port 1: presure.");
        for (i_stimulus_port1 = 0; i_stimulus_port1 < 100; i_stimulus_port1 = i_stimulus_port1 + 1) begin
            $display ("Port 1 Send: 3->2 #0d ", i_stimulus_port1);
            if (mac_speed[1] == 2'b10) begin
                send_frame_1g_port1(frame2.tobits(0), i_stimulus_port1);
            end
            else if(mac_speed[1] == 2'b01) begin
                send_frame_100m_port1(frame2.tobits(0), i_stimulus_port1);
            end

        end

        // wait (tx_monitor_finished_1G == 4'b1111);
        rx_stimulus_pressure_finished[1] = 1;
        #10;
    end // p_rx_stimulus_port1

    integer i_stimulus_port2;

    initial
    begin : p_rx_stimulus_port2
        wait(rx_stimulus_warmup_finished == 1);
        #10;

        // 1 Gb/s speed
        //-----------------------------------------------------
        
        // Presure test
        $display("Phase two of stimulation port 2: presure.");
        for (i_stimulus_port2 = 0; i_stimulus_port2 < 100; i_stimulus_port2 = i_stimulus_port2 + 1) begin
            $display ("Port 2 Send: 2->1 #0d ", i_stimulus_port2);
            if (mac_speed[2] == 2'b10) begin
                send_frame_1g_port2(frame1.tobits(0), i_stimulus_port2);
            end
            else if(mac_speed[2] == 2'b01) begin
                send_frame_100m_port2(frame1.tobits(0), i_stimulus_port2);
            end

        end

        // wait (tx_monitor_finished_1G == 4'b1111);
        rx_stimulus_pressure_finished[2] = 1;
        #10;
    end // p_rx_stimulus_port2

    integer i_stimulus_port3;

    initial
    begin : p_rx_stimulus_port3
        wait(rx_stimulus_warmup_finished == 1);
        #10;

        // 1 Gb/s speed
        //-----------------------------------------------------

        // Presure test
        // $display("Phase two of stimulation port 3: presure.");
        // for (i_stimulus_port3 = 0; i_stimulus_port3 < 100; i_stimulus_port3 = i_stimulus_port3 + 1) begin
        //     $display ("Send 3->0:#0d ", i_stimulus_port3);
        //     if (mac_speed[3] == 2'b10) begin
        //         send_frame_1g_port3(frame1.tobits(0), i_stimulus_port3);
        //     end
        //     else if(mac_speed[3] == 2'b01) begin
        //         send_frame_100m_port3(frame1.tobits(0), i_stimulus_port3);
        //     end
        // end

        // wait (tx_monitor_finished_1G == 4'b1111);
        rx_stimulus_pressure_finished[3] = 1;
        #10;
    end // p_rx_stimulus


    //----------------------------------------------------------------------------
    // A Task to check a transmitted frame at 1Gb/s
    //----------------------------------------------------------------------------
    task check_frame_1g_port0;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[0] !== 1'b1)
            @(rgmii_txc[0]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[0]) begin
            $display("** ERROR: tx_ctl[0] started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[0] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[0] === 4'h5)
            @(negedge rgmii_txc[0]);

        // Parse over the SFD
        if (rgmii_txd[0] !== 4'hd) begin
            $display("** ERROR: Port 0, SFD not present at %t", $realtime, "ps");
            demo_mode_error[0] <= 1;
        end
        @(posedge rgmii_txc[0]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[0][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[0];
                @(rgmii_txc[0]);
                rgmii_column[7:4] = rgmii_txd[0][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[0];
                
                tx_monitor_working_frame_0.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_0.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_0.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[0]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_0.data[12];
            frame_length[7:0] = tx_monitor_working_frame_0.data[13];

            // while (column_index <  frame_length + 14) begin
            while (rgmii_tx_ctl[0] == 1'b1) begin
                rgmii_column[3:0] = rgmii_txd[0][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[0];
                @(rgmii_txc[0]);
                rgmii_column[7:4] = rgmii_txd[0][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[0];
                
                tx_monitor_working_frame_0.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_0.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_0.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[0]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            for (I = 0; I < 4; I = I + 1)
            begin
                rgmii_column[3:0] = rgmii_txd[0][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[0];
                @(rgmii_txc[0]);
                rgmii_column[7:4] = rgmii_txd[0][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[0];

                if (rgmii_valid !== 2'b11) begin
                    $display("** ERROR: rgmii_tx_ctl[0] incorrect during FCS field at %t", $realtime, "ps");
                    demo_mode_error[0] <= 1;
                end

                case(I)
                    0 : if (rgmii_column !== fcs[7:0]) begin
                            $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[0] <= 1;
                        end
                    1 :  if (rgmii_column !== fcs[15:8]) begin
                            $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[0] <= 1;
                        end
                    2 :  if (rgmii_column !== fcs[23:16]) begin
                            $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[0] <= 1;
                        end
                    3 :  if (rgmii_column !== fcs[31:24]) begin
                            $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[0] <= 1;
                        end
                endcase
                @(rgmii_txc[0]);
            end

            dst_mac[47:40] = tx_monitor_working_frame_0.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_0.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_0.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_0.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_0.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_0.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_0.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_0.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_0.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_0.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_0.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_0.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_0.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_0.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_0.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_0.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 0 recv packet.\nDst mac: %h, Src mac: %h.\nSeq:%h.", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_1g_port0

    task check_frame_1g_port1;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[1] !== 1'b1)
            @(rgmii_txc[1]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[1]) begin
            $display("** ERROR: tx_ctl[1] started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[1] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[1] === 4'h5)
            @(negedge rgmii_txc[1]);

        // Parse over the SFD
        if (rgmii_txd[1] !== 4'hd) begin
            $display("** ERROR: Port 1, SFD not present at %t", $realtime, "ps");
            demo_mode_error[1] <= 1;
        end
        @(posedge rgmii_txc[1]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[1][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[1];
                @(rgmii_txc[1]);
                rgmii_column[7:4] = rgmii_txd[1][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[1];
                
                tx_monitor_working_frame_1.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_1.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_1.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[1]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_1.data[12];
            frame_length[7:0] = tx_monitor_working_frame_1.data[13];

            while (column_index <  frame_length + 14) begin
                rgmii_column[3:0] = rgmii_txd[1][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[1];
                @(rgmii_txc[1]);
                rgmii_column[7:4] = rgmii_txd[1][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[1];
                
                tx_monitor_working_frame_1.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_1.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_1.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[1]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            for (I = 0; I < 4; I = I + 1)
            begin
                rgmii_column[3:0] = rgmii_txd[1][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[1];
                @(rgmii_txc[1]);
                rgmii_column[7:4] = rgmii_txd[1][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[1];

                if (rgmii_valid !== 2'b11) begin
                    $display("** ERROR: rgmii_tx_ctl[1] incorrect during FCS field at %t", $realtime, "ps");
                    demo_mode_error[1] <= 1;
                end

                case(I)
                    0 : if (rgmii_column !== fcs[7:0]) begin
                            $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[1] <= 1;
                        end
                    1 :  if (rgmii_column !== fcs[15:8]) begin
                            $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[1] <= 1;
                        end
                    2 :  if (rgmii_column !== fcs[23:16]) begin
                            $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[1] <= 1;
                        end
                    3 :  if (rgmii_column !== fcs[31:24]) begin
                            $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[1] <= 1;
                        end
                endcase
                @(rgmii_txc[1]);
            end

            dst_mac[47:40] = tx_monitor_working_frame_1.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_1.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_1.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_1.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_1.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_1.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_1.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_1.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_1.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_1.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_1.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_1.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_1.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_1.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_1.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_1.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 1 recv packet.\nDst mac: %h, Src mac: %h.\nSeq:%h.", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_1g_port1

    task check_frame_1g_port2;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[2] !== 1'b1)
            @(rgmii_txc[2]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[2]) begin
            $display("** ERROR: tx_ctl[2] started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[2] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[2] === 4'h5)
            @(negedge rgmii_txc[2]);

        // Parse over the SFD
        if (rgmii_txd[2] !== 4'hd) begin
            $display("** ERROR: Port 2, SFD not present at %t", $realtime, "ps");
            demo_mode_error[2] <= 1;
        end
        @(posedge rgmii_txc[2]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[2][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[2];
                @(rgmii_txc[2]);
                rgmii_column[7:4] = rgmii_txd[2][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[2];
                
                tx_monitor_working_frame_2.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_2.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_2.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[2]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_2.data[12];
            frame_length[7:0] = tx_monitor_working_frame_2.data[13];

            while (column_index <  frame_length + 14) begin
                rgmii_column[3:0] = rgmii_txd[2][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[2];
                @(rgmii_txc[2]);
                rgmii_column[7:4] = rgmii_txd[2][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[2];
                
                tx_monitor_working_frame_2.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_2.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_2.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[2]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            for (I = 0; I < 4; I = I + 1)
            begin
                rgmii_column[3:0] = rgmii_txd[2][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[2];
                @(rgmii_txc[2]);
                rgmii_column[7:4] = rgmii_txd[2][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[2];

                if (rgmii_valid !== 2'b11) begin
                    $display("** ERROR: rgmii_tx_ctl[2] incorrect during FCS field at %t", $realtime, "ps");
                    demo_mode_error[2] <= 1;
                end

                case(I)
                    0 : if (rgmii_column !== fcs[7:0]) begin
                            $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[2] <= 1;
                        end
                    1 :  if (rgmii_column !== fcs[15:8]) begin
                            $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[2] <= 1;
                        end
                    2 :  if (rgmii_column !== fcs[23:16]) begin
                            $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[2] <= 1;
                        end
                    3 :  if (rgmii_column !== fcs[31:24]) begin
                            $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[2] <= 1;
                        end
                endcase
                @(rgmii_txc[2]);
            end

            dst_mac[47:40] = tx_monitor_working_frame_2.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_2.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_2.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_2.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_2.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_2.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_2.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_2.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_2.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_2.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_2.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_2.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_2.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_2.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_2.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_2.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 2 recv packet.\nDst mac: %h, Src mac: %h.\nSeq:%h.", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_1g_port2

    task check_frame_1g_port3;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[3] !== 1'b1)
            @(rgmii_txc[3]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[3]) begin
            $display("** ERROR: tx_ctl[3] started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[3] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[3] === 4'h5)
            @(negedge rgmii_txc[3]);

        // Parse over the SFD
        if (rgmii_txd[3] !== 4'hd) begin
            $display("** ERROR: Port 3, SFD not present at %t", $realtime, "ps");
            demo_mode_error[3] <= 1;
        end
        @(posedge rgmii_txc[3]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[3][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[3];
                @(rgmii_txc[3]);
                rgmii_column[7:4] = rgmii_txd[3][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[3];
                
                tx_monitor_working_frame_3.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_3.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_3.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[3]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_3.data[12];
            frame_length[7:0] = tx_monitor_working_frame_3.data[13];

            while (column_index <  frame_length + 14) begin
                rgmii_column[3:0] = rgmii_txd[3][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[3];
                @(rgmii_txc[3]);
                rgmii_column[7:4] = rgmii_txd[3][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[3];
                
                tx_monitor_working_frame_3.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_3.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_3.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(rgmii_txc[3]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            for (I = 0; I < 4; I = I + 1)
            begin
                rgmii_column[3:0] = rgmii_txd[3][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[3];
                @(rgmii_txc[3]);
                rgmii_column[7:4] = rgmii_txd[3][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[3];

                if (rgmii_valid !== 2'b11) begin
                    $display("** ERROR: rgmii_tx_ctl[3] incorrect during FCS field at %t", $realtime, "ps");
                    demo_mode_error[3] <= 1;
                end

                case(I)
                    0 : if (rgmii_column !== fcs[7:0]) begin
                            $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[3] <= 1;
                        end
                    1 :  if (rgmii_column !== fcs[15:8]) begin
                            $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[3] <= 1;
                        end
                    2 :  if (rgmii_column !== fcs[23:16]) begin
                            $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[3] <= 1;
                        end
                    3 :  if (rgmii_column !== fcs[31:24]) begin
                            $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
                            demo_mode_error[3] <= 1;
                        end
                endcase
                @(rgmii_txc[3]);
            end

            dst_mac[47:40] = tx_monitor_working_frame_3.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_3.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_3.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_3.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_3.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_3.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_3.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_3.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_3.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_3.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_3.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_3.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_3.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_3.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_3.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_3.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 3 recv packet.\nDst mac: %h, Src mac: %h.\nSeq:%h.", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_1g_port3

    //----------------------------------------------------------------------------
    // A Task to check a transmitted frame at 1Gb/s
    //----------------------------------------------------------------------------
    task check_frame_100m_port0;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[0] !== 1'b1)
            @(posedge rgmii_txc[0]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[0]) begin
            $display("** ERROR: tx_ctl started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[0] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[0] === 4'h5)
            @(negedge rgmii_txc[0]);

        // Parse over the SFD
        if (rgmii_txd[0] !== 4'hd) begin
            $display("** ERROR: Port 0, SFD not present at %t", $realtime, "ps");
            demo_mode_error[0] <= 1;
        end
        @(posedge rgmii_txc[0]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[0][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[0];
                @(posedge rgmii_txc[0]);
                rgmii_column[7:4] = rgmii_txd[0][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[0];
                
                tx_monitor_working_frame_0.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_0.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_0.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[0]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_0.data[12];
            frame_length[7:0] = tx_monitor_working_frame_0.data[13];

            // while (column_index <  frame_length + 14) begin
            while (rgmii_tx_ctl[0] == 1'b1) begin
                rgmii_column[3:0] = rgmii_txd[0][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[0];
                @(posedge rgmii_txc[0]);
                rgmii_column[7:4] = rgmii_txd[0][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[0];
                
                tx_monitor_working_frame_0.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_0.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_0.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[0]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            // for (I = 0; I < 4; I = I + 1)
            // begin
            //     rgmii_column[3:0] = rgmii_txd[0][3:0];
            //     rgmii_valid[0]    = rgmii_tx_ctl[0];
            //     @(posedge rgmii_txc[0]);
            //     rgmii_column[7:4] = rgmii_txd[0][3:0];
            //     rgmii_valid[1]    = rgmii_tx_ctl[0];

            //     if (rgmii_valid !== 2'b11) begin
            //         $display("** ERROR: rgmii_tx_ctl[0] incorrect during FCS field at %t", $realtime, "ps");
            //         demo_mode_error[0] <= 1;
            //     end

            //     case(I)
            //         0 : if (rgmii_column !== fcs[7:0]) begin
            //                 $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[0] <= 1;
            //             end
            //         1 :  if (rgmii_column !== fcs[15:8]) begin
            //                 $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[0] <= 1;
            //             end
            //         2 :  if (rgmii_column !== fcs[23:16]) begin
            //                 $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[0] <= 1;
            //             end
            //         3 :  if (rgmii_column !== fcs[31:24]) begin
            //                 $display("** ERROR: rgmii_txd[0] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[0] <= 1;
            //             end
            //     endcase
            //     @(posedge rgmii_txc[0]);
            // end

            dst_mac[47:40] = tx_monitor_working_frame_0.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_0.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_0.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_0.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_0.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_0.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_0.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_0.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_0.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_0.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_0.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_0.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_0.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_0.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_0.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_0.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, " Port 0 recv packet.\nDst mac: %h, Src mac: %h.\n", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_100m_port0

    task check_frame_100m_port1;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[1] !== 1'b1)
            @(posedge rgmii_txc[1]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[1]) begin
            $display("** ERROR: tx_ctl started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[1] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[1] === 4'h5)
            @(negedge rgmii_txc[1]);

        // Parse over the SFD
        if (rgmii_txd[1] !== 4'hd) begin
            $display("** ERROR: Port 0, SFD not present at %t", $realtime, "ps");
            demo_mode_error[1] <= 1;
        end
        @(posedge rgmii_txc[1]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[1][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[1];
                @(posedge rgmii_txc[1]);
                rgmii_column[7:4] = rgmii_txd[1][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[1];
                
                tx_monitor_working_frame_1.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_1.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_1.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[1]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_1.data[12];
            frame_length[7:0] = tx_monitor_working_frame_1.data[13];

            // while (column_index <  frame_length + 14) begin
            while (rgmii_tx_ctl[1] == 1'b1) begin
                // if (rgmii_tx_ctl[1] != 1'b1) begin
                //     break;
                // end
                rgmii_column[3:0] = rgmii_txd[1][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[1];
                @(posedge rgmii_txc[1]);
                rgmii_column[7:4] = rgmii_txd[1][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[1];
                
                tx_monitor_working_frame_1.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_1.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_1.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[1]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            // for (I = 0; I < 4; I = I + 1)
            // begin
            //     rgmii_column[3:0] = rgmii_txd[1][3:0];
            //     rgmii_valid[0]    = rgmii_tx_ctl[1];
            //     @(posedge rgmii_txc[1]);
            //     rgmii_column[7:4] = rgmii_txd[1][3:0];
            //     rgmii_valid[1]    = rgmii_tx_ctl[1];

            //     if (rgmii_valid !== 2'b11) begin
            //         $display("** ERROR: rgmii_tx_ctl[1] incorrect during FCS field at %t", $realtime, "ps");
            //         demo_mode_error[1] <= 1;
            //     end

            //     case(I)
            //         0 : if (rgmii_column !== fcs[7:0]) begin
            //                 $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[1] <= 1;
            //             end
            //         1 :  if (rgmii_column !== fcs[15:8]) begin
            //                 $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[1] <= 1;
            //             end
            //         2 :  if (rgmii_column !== fcs[23:16]) begin
            //                 $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[1] <= 1;
            //             end
            //         3 :  if (rgmii_column !== fcs[31:24]) begin
            //                 $display("** ERROR: rgmii_txd[1] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[1] <= 1;
            //             end
            //     endcase
            //     @(posedge rgmii_txc[1]);
            // end

            dst_mac[47:40] = tx_monitor_working_frame_1.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_1.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_1.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_1.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_1.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_1.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_1.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_1.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_1.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_1.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_1.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_1.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_1.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_1.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_1.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_1.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 1 recv packet.\nDst mac: %h, Src mac: %h.\nSeq:%h.", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_100m_port1

    task check_frame_100m_port2;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[2] !== 1'b1)
            @(posedge rgmii_txc[2]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[2]) begin
            $display("** ERROR: tx_ctl started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[2] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[2] === 4'h5)
            @(negedge rgmii_txc[2]);

        // Parse over the SFD
        if (rgmii_txd[2] !== 4'hd) begin
            $display("** ERROR: Port 0, SFD not present at %t", $realtime, "ps");
            demo_mode_error[2] <= 1;
        end
        @(posedge rgmii_txc[2]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[2][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[2];
                @(posedge rgmii_txc[2]);
                rgmii_column[7:4] = rgmii_txd[2][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[2];
                
                tx_monitor_working_frame_2.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_2.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_2.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[2]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_2.data[12];
            frame_length[7:0] = tx_monitor_working_frame_2.data[13];

            // while (column_index <  frame_length + 14) begin
            while (rgmii_tx_ctl[2] == 1'b1) begin
                // if (rgmii_tx_ctl[2] != 1'b1) begin
                //     break;
                // end
                rgmii_column[3:0] = rgmii_txd[2][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[2];
                @(posedge rgmii_txc[2]);
                rgmii_column[7:4] = rgmii_txd[2][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[2];
                
                tx_monitor_working_frame_2.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_2.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_2.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[2]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            // for (I = 0; I < 4; I = I + 1)
            // begin
            //     rgmii_column[3:0] = rgmii_txd[2][3:0];
            //     rgmii_valid[0]    = rgmii_tx_ctl[2];
            //     @(posedge rgmii_txc[2]);
            //     rgmii_column[7:4] = rgmii_txd[2][3:0];
            //     rgmii_valid[1]    = rgmii_tx_ctl[2];

            //     if (rgmii_valid !== 2'b11) begin
            //         $display("** ERROR: rgmii_tx_ctl[2] incorrect during FCS field at %t", $realtime, "ps");
            //         demo_mode_error[2] <= 1;
            //     end

            //     case(I)
            //         0 : if (rgmii_column !== fcs[7:0]) begin
            //                 $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[2] <= 1;
            //             end
            //         1 :  if (rgmii_column !== fcs[15:8]) begin
            //                 $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[2] <= 1;
            //             end
            //         2 :  if (rgmii_column !== fcs[23:16]) begin
            //                 $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[2] <= 1;
            //             end
            //         3 :  if (rgmii_column !== fcs[31:24]) begin
            //                 $display("** ERROR: rgmii_txd[2] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[2] <= 1;
            //             end
            //     endcase
            //     @(posedge rgmii_txc[2]);
            // end

            dst_mac[47:40] = tx_monitor_working_frame_2.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_2.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_2.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_2.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_2.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_2.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_2.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_2.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_2.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_2.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_2.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_2.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_2.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_2.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_2.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_2.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 2 recv packet.\nDst mac: %h, Src mac: %h.\n", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_100m_port2

    task check_frame_100m_port3;
        integer column_index;
        integer I;
        integer frame_length;
        reg [31:0] fcs;
        reg [7:0]  rgmii_column;
        reg [1:0]  rgmii_valid;
        reg [47:0] dst_mac;
        reg [47:0] src_mac;
        reg [31:0] seq_num;
    begin
        column_index = 0;
        frame_length = 0;

        // reset the fcs calculation
        fcs = 32'b0;

        // wait until the first real column of data to come out of RX client
        while (rgmii_tx_ctl[3] !== 1'b1)
            @(posedge rgmii_txc[3]);

        // check tx_ctl has gone high at the correct edge (should be rising)
        if (!rgmii_txc[3]) begin
            $display("** ERROR: tx_ctl started on incorrect phase at %t", $realtime, "ps");
            demo_mode_error[3] <= 1;
        end

        // Parse over the preamble field
        while (rgmii_txd[3] === 4'h5)
            @(negedge rgmii_txc[3]);

        // Parse over the SFD
        if (rgmii_txd[3] !== 4'hd) begin
            $display("** ERROR: Port 0, SFD not present at %t", $realtime, "ps");
            demo_mode_error[3] <= 1;
        end
        @(posedge rgmii_txc[3]);

        if (TB_MODE == "DEMO") begin
            // Receive Ethernet header
            while (column_index < 14) begin
                rgmii_column[3:0] = rgmii_txd[3][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[3];
                @(posedge rgmii_txc[3]);
                rgmii_column[7:4] = rgmii_txd[3][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[3];
                
                tx_monitor_working_frame_3.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_3.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_3.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[3]);
            end

            // Receive following data based on Length field.
            frame_length[15:8] = tx_monitor_working_frame_3.data[12];
            frame_length[7:0] = tx_monitor_working_frame_3.data[13];

            // while (column_index <  frame_length + 14) begin
            // while (1'b1) begin
            while (rgmii_tx_ctl[3] == 1'b1) begin
                rgmii_column[3:0] = rgmii_txd[3][3:0];
                rgmii_valid[0]    = rgmii_tx_ctl[3];
                @(posedge rgmii_txc[3]);
                rgmii_column[7:4] = rgmii_txd[3][3:0];
                rgmii_valid[1]    = rgmii_tx_ctl[3];
                
                tx_monitor_working_frame_3.valid[column_index] = rgmii_valid[0];
                tx_monitor_working_frame_3.error[column_index] = rgmii_valid[1] ^ rgmii_valid[0];
                tx_monitor_working_frame_3.data[column_index] = rgmii_column;

                // calculate expected crc for the frame
                calc_crc(rgmii_column, fcs);

                // wait for next column of data
                column_index = column_index + 1;
                @(posedge rgmii_txc[3]);
            end

            // Check the FCS
            // Having checked all data columns, txd must contain FCS.
            // for (I = 0; I < 4; I = I + 1)
            // begin
            //     rgmii_column[3:0] = rgmii_txd[3][3:0];
            //     rgmii_valid[0]    = rgmii_tx_ctl[3];
            //     @(posedge rgmii_txc[3]);
            //     rgmii_column[7:4] = rgmii_txd[3][3:0];
            //     rgmii_valid[1]    = rgmii_tx_ctl[3];

            //     if (rgmii_valid !== 2'b11) begin
            //         $display("** ERROR: rgmii_tx_ctl[3] incorrect during FCS field at %t", $realtime, "ps");
            //         demo_mode_error[3] <= 1;
            //     end

            //     case(I)
            //         0 : if (rgmii_column !== fcs[7:0]) begin
            //                 $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[3] <= 1;
            //             end
            //         1 :  if (rgmii_column !== fcs[15:8]) begin
            //                 $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[3] <= 1;
            //             end
            //         2 :  if (rgmii_column !== fcs[23:16]) begin
            //                 $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[3] <= 1;
            //             end
            //         3 :  if (rgmii_column !== fcs[31:24]) begin
            //                 $display("** ERROR: rgmii_txd[3] incorrect during FCS field at %t", $realtime, "ps");
            //                 demo_mode_error[3] <= 1;
            //             end
            //     endcase
            //     @(posedge rgmii_txc[3]);
            // end

            dst_mac[47:40] = tx_monitor_working_frame_3.data[0][7:0];
            dst_mac[39:32] = tx_monitor_working_frame_3.data[1][7:0];
            dst_mac[31:24] = tx_monitor_working_frame_3.data[2][7:0];
            dst_mac[23:16] = tx_monitor_working_frame_3.data[3][7:0];
            dst_mac[15:8] = tx_monitor_working_frame_3.data[4][7:0];
            dst_mac[7:0] = tx_monitor_working_frame_3.data[5][7:0];

            src_mac[47:40] = tx_monitor_working_frame_3.data[6][7:0];
            src_mac[39:32] = tx_monitor_working_frame_3.data[7][7:0];
            src_mac[31:24] = tx_monitor_working_frame_3.data[8][7:0];
            src_mac[23:16] = tx_monitor_working_frame_3.data[9][7:0];
            src_mac[15:8] = tx_monitor_working_frame_3.data[10][7:0];
            src_mac[7:0] = tx_monitor_working_frame_3.data[11][7:0];

            seq_num[31:24] = tx_monitor_working_frame_3.data[SEQ_OFFSET];
            seq_num[23:16] = tx_monitor_working_frame_3.data[SEQ_OFFSET+1];
            seq_num[15:8] = tx_monitor_working_frame_3.data[SEQ_OFFSET+2];
            seq_num[7:0] = tx_monitor_working_frame_3.data[SEQ_OFFSET+3];
            // Have received the frame. Now print useful information.
            $display($time, "Port 3 recv packet.\nDst mac: %h, Src mac: %h.\n", dst_mac, src_mac, seq_num);
        end
    end
    endtask // check_frame_100m_port3

    //----------------------------------------------------------------------------
    // Monitor process. This process checks the data coming out of the
    // transmitter to make sure that it matches that inserted into the
    // receiver.
    //----------------------------------------------------------------------------

    // Monitor process for port 0
    initial
    begin : p_tx_monitor_0
        // wait for the reset to complete before starting monitor
        @(negedge reset);

        // Check the frames
        while (1) begin
            if (mac_speed[0] == 2'b10) begin
                check_frame_1g_port0();
            end
            else if (mac_speed[0] == 2'b01) begin
                check_frame_100m_port0();
            end
        end
    end // p_tx_monitor_port0

    // Monitor process for port 1
    initial
    begin : p_tx_monitor_1
        // wait for the reset to complete before starting monitor
        @(negedge reset);

        // Check the frames
        while (1) begin
            if (mac_speed[0] == 2'b10) begin
                check_frame_1g_port1();
            end
            else if (mac_speed[0] == 2'b01) begin
                check_frame_100m_port1();
            end
        end
    end // p_tx_monitor_port1

    // Monitor process for port 2
    initial
    begin : p_tx_monitor_2
        // wait for the reset to complete before starting monitor
        @(negedge reset);

        // Check the frames
        while (1) begin
            if (mac_speed[0] == 2'b10) begin
                check_frame_1g_port2();
            end
            else if (mac_speed[0] == 2'b01) begin
                check_frame_100m_port2();
            end
        end
    end // p_tx_monitor_port2

    // Monitor process for port 3
    initial
    begin : p_tx_monitor_3
        // wait for the reset to complete before starting monitor
        @(negedge reset);

        // Check the frames
        while (1) begin
            if (mac_speed[0] == 2'b10) begin
                check_frame_1g_port3();
            end
            else if (mac_speed[0] == 2'b01) begin
                check_frame_100m_port3();
            end
        end
    end // p_tx_monitor_port3

    // parameter integer C_M_AXI_ADDR_WIDTH = 32;
    // parameter integer C_M_AXI_DATA_WIDTH = 32;

    // // System Signals
    // wire M_AXI_ACLK;
    // wire M_AXI_ARESETN;

    // // Master Interface Write Address
    // wire [C_M_AXI_ADDR_WIDTH-1:0] M_AXI_AWADDR;
    // wire [3-1:0] M_AXI_AWPROT;
    // wire M_AXI_AWVALID;
    // wire M_AXI_AWREADY;

    // // Master Interface Write Data
    // wire [C_M_AXI_DATA_WIDTH-1:0] M_AXI_WDATA;
    // wire [C_M_AXI_DATA_WIDTH/8-1:0] M_AXI_WSTRB;
    // wire M_AXI_WVALID;
    // wire M_AXI_WREADY;

    // // Master Interface Write Response
    // wire [2-1:0] M_AXI_BRESP;
    // wire M_AXI_BVALID;
    // wire M_AXI_BREADY;

    // // Master Interface Read Address
    // wire [C_M_AXI_ADDR_WIDTH-1:0] M_AXI_ARADDR;
    // wire [3-1:0] M_AXI_ARPROT;
    // wire M_AXI_ARVALID;
    // wire M_AXI_ARREADY;

    // // Master Interface Read Data 
    // wire [C_M_AXI_DATA_WIDTH-1:0] M_AXI_RDATA;
    // wire [2-1:0] M_AXI_RRESP;
    // wire M_AXI_RVALID;
    // wire M_AXI_RREADY;

    // // External Signals
    // wire INTR_IN;

    // // AXI4 signals
    // reg 		awvalid;
    // reg 		wvalid;
    // reg 		push_write;
    // reg 		pop_read;
    // reg          arvalid;
    // reg          rready;
    // reg          bready;
    // reg [31:0] 	awaddr;
    // reg [31:0] 	wdata;
    // reg [31:0] 	araddr;
    // wire 	write_resp_error;
    // wire         read_resp_error;
    
    // /////////////////
    // //I/O Connections
    // /////////////////
    // //////////////////// 
    // //Write Address (AW)
    // ////////////////////
    // assign M_AXI_AWADDR = awaddr;
    
    // assign M_AXI_WDATA = wdata;
    // assign M_AXI_AWPROT = 3'h0;
    // assign M_AXI_AWVALID = awvalid;

    // ///////////////
    // //Write Data(W)
    // ///////////////
    // assign M_AXI_WVALID = wvalid;

    // //Set all byte strobes in this example
    // assign M_AXI_WSTRB = -1;

    // ////////////////////
    // //Write Response (B)
    // ////////////////////
    // assign M_AXI_BREADY = bready;

    // ///////////////////   
    // //Read Address (AR)
    // ///////////////////
    // assign M_AXI_ARADDR = araddr;
    // assign M_AXI_ARVALID = arvalid;
    // assign M_AXI_ARPROT = 3'b0;

    // ////////////////////////////
    // //Read and Read Response (R)
    // ////////////////////////////
    // assign M_AXI_RREADY = rready;
    
    // ///////////////////////
    // //Write Address Channel
    // ///////////////////////
    // /*
    // The purpose of the write address channel is to request the address and 
    // command information for the entire transaction.  It is a single beat
    // of information.
    
    // Note for this example the awvalid/wvalid are asserted at the same
    // time, and then each is deasserted independent from each other.
    // This is a lower-performance, but simplier control scheme.
    
    // AXI VALID signals must be held active until accepted by the partner.
    
    // A data transfer is accepted by the slave when a master has
    // VALID data and the slave acknoledges it is also READY. While the master
    // is allowed to generated multiple, back-to-back requests by not 
    // deasserting VALID, this design will add an extra rest cycle for
    // simplicity.
    
    // Since only one outstanding transaction is issued by the user design,
    // there will not be a collision between a new request and an accepted
    // request on the same clock cycle. Otherwise, an additional clause is 
    // necessary.
    // */
    // always @(posedge M_AXI_ACLK)
    // begin
        
    //     //Only VALID signals must be deasserted during reset per AXI spec
    //     //Consider inverting then registering active-low reset for higher fmax
    //     if (M_AXI_ARESETN == 0 )
    //     awvalid <= 1'b0;

    //     //Address accepted by interconnect/slave
    //     else if (M_AXI_AWREADY && awvalid)
    //     awvalid <= 1'b0;

    //     //Signal a new address/data command is available by user logic
    //     else if (push_write)
    //     awvalid <= 1'b1;
    //     else
    //     awvalid <= awvalid;
    // end 

    // ////////////////////
    // //Write Data Channel
    // ////////////////////
    // /*
    // The write data channel is for transfering the actual data.
    
    // The data generation is specific to the example design, and
    // so only the WVALID/WREADY handshake is shown here
    // */
    // always @(posedge M_AXI_ACLK)
    // begin
    //     if (M_AXI_ARESETN == 0 )
    //     wvalid <= 1'b0;
        
    //     //Data accepted by interconnect/slave
    //     else if (M_AXI_WREADY && wvalid)
    //     wvalid <= 1'b0;

    //     //Signal a new address/data command is available by user logic
    //     else if (push_write)
    //     wvalid <= 1'b1;
    //     else
    //     wvalid <= awvalid;
    // end 

    // ////////////////////////////
    // //Write Response (B) Channel
    // ////////////////////////////
    // /* 
    // The write response channel provides feedback that the write has committed
    // to memory. BREADY will occur after both the data and the write address
    // has arrived and been accepted by the slave, and can guarantee that no
    // other accesses launched afterwards will be able to be reordered before it.
    
    // The BRESP bit [1] is used indicate any errors from the interconnect or
    // slave for the entire write burst. This example will capture the error.
    
    // While not necessary per spec, it is advisable to reset READY signals in
    // case of differing reset latencies between master/slave.
    // */

    // //Always accept write responses
    // always @(posedge M_AXI_ACLK)
    // begin
    //     if (M_AXI_ARESETN == 0)
    //     bready <= 1'b0;
    //     else
    //     bready <= 1'b1;
    // end

    // //Flag write errors
    // assign write_resp_error = bready & M_AXI_BVALID & M_AXI_BRESP[1];
    
    // //////////////////////   
    // //Read Address Channel
    // //////////////////////
    // always @(posedge M_AXI_ACLK)
    // begin
    //     if (M_AXI_ARESETN == 0 )
    //     arvalid <= 1'b0;
    //     else if (M_AXI_ARREADY && arvalid)
    //     arvalid <= 1'b0;
    //     else if (pop_read)
    //     arvalid <= 1'b1;
    //     else
    //     arvalid <= arvalid;
    // end 

    // //////////////////////////////////   
    // //Read Data (and Response) Channel
    // //////////////////////////////////
    // /* 
    // The Read Data channel returns the results of the read request 
    
    // In this example the data checker is always able to accept
    // more data, so no need to throttle the RREADY signal. 
    
    // While not necessary per spec, it is advisable to reset READY signals in
    // case of differing reset latencies between master/slave.
    // */ 
    // always @(posedge M_AXI_ACLK)
    // begin
    //     if (M_AXI_ARESETN == 0)
    //     rready <= 1'b0;
    //     else
    //     rready <= 1'b1;
    // end

    // //Flag write errors
    // assign read_resp_error = rready & M_AXI_RVALID & M_AXI_RRESP[1];  

    // ////////////
    // //User Logic
    // ////////////

    // ///////////////////////
    // //Main write controller
    // ///////////////////////
    // /*  
    // By only issuing one request at a time, the control logic is 
    // simplified.
    
    // Request a new write if:
    // -A command was not just submitted
    // -AW and W channels are both idle
    // -A new request was not requested last cycle
    // */
    // /*always @(posedge M_AXI_ACLK)
    // begin
    //     if (M_AXI_ARESETN == 0 )
    //     begin
    //     push_write <= 1'b0;
    //     end

    //     //Request new write
    //     else if (~awvalid && ~wvalid && ~push_write)
    //     begin
    //     push_write <= 1'b1;
    //     end
    //     else
    //     begin
    //     push_write <= 1'b0; //Negate to generate a pulse
    //     end
    // end */

    // //////////////////////
    // //Main read controller
    // //////////////////////
    // /*
    // By only issuing one request at a time, the control logic is 
    // simplified.

    // Request a new read if:
    // -A command was not just submitted
    // -AR channel is idle
    // -A new request was not requested last cycle
    // */
    // /*always @(posedge M_AXI_ACLK)
    // begin
    //     if (M_AXI_ARESETN == 0 )
    //     begin
    //     pop_read <= 1'b0;
    //     end

    //     //Request new read
    //     else if (~arvalid && ~pop_read)
    //     begin
    //     pop_read <= 1'b1;	  
    //     end
    //     else
    //     begin
    //     pop_read <= 1'b0; //Negate to generate a pulse
    //     end
    // end */


    // task axi4_wr_req(input [31:0]addr, input [31:0]data);
    // integer i;
    // begin
    // $write("axi4_wr %08x", addr);
    // $write(" %08x", data);
    // for (i=0; i<1; i=i+1) @(posedge M_AXI_ACLK);
    // awaddr     = addr;
    // wdata      = data;
    // push_write = 1'b1;
    // for (i=0; i<1; i=i+1) @(posedge M_AXI_ACLK);
    // awaddr     = addr;
    // wdata      = data;
    // push_write = 1'b0;
    // for (i=0; i<1; i=i+1) @(posedge M_AXI_ACLK);
    // @(~awvalid && ~wvalid);
    // end
    // endtask

    // task axi4_rd_req(input [31:0]addr);
    // integer i;
    // begin
    // $write("axi4_rd %08x", addr);
    // for (i=0; i<1; i=i+1) @(posedge M_AXI_ACLK);
    // araddr   = addr;
    // pop_read = 1'b1;
    // for (i=0; i<1; i=i+1) @(posedge M_AXI_ACLK);
    // araddr   = addr;
    // pop_read = 1'b0;
    // for (i=0; i<1; i=i+1) @(posedge M_AXI_ACLK);
    // @(~arvalid);
    // end
    // endtask

    // task axi4_wr_ack;
    // begin
    // @(M_AXI_BVALID && bready);
    // @(posedge M_AXI_ACLK);
    // $write(" W_RESP: %08x\n", M_AXI_BRESP);
    // end
    // endtask

    // task axi4_rd_ack;
    // begin
    // @(M_AXI_RVALID && rready);
    // @(posedge M_AXI_ACLK);
    // $write(" %08x", M_AXI_RDATA);
    // $write(" R_RESP: %08x\n", M_AXI_RRESP);
    // end
    // endtask

    // initial begin
    // #300;
    // @(posedge M_AXI_ACLK);
    // axi4_wr_req(32'h00000004,32'h12345678);axi4_wr_ack;
    // axi4_rd_req(32'h00000004             );axi4_rd_ack;
    // end
endmodule
